VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fibonacci
  CLASS BLOCK ;
  FOREIGN fibonacci ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.280 0.000 763.840 4.000 ;
    END
  END clk
  PIN fn[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 596.000 16.240 600.000 ;
    END
  END fn[0]
  PIN fn[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 596.000 296.240 600.000 ;
    END
  END fn[10]
  PIN fn[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 596.000 324.240 600.000 ;
    END
  END fn[11]
  PIN fn[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 596.000 352.240 600.000 ;
    END
  END fn[12]
  PIN fn[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 596.000 380.240 600.000 ;
    END
  END fn[13]
  PIN fn[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 596.000 408.240 600.000 ;
    END
  END fn[14]
  PIN fn[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 596.000 436.240 600.000 ;
    END
  END fn[15]
  PIN fn[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 596.000 464.240 600.000 ;
    END
  END fn[16]
  PIN fn[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 596.000 492.240 600.000 ;
    END
  END fn[17]
  PIN fn[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 519.680 596.000 520.240 600.000 ;
    END
  END fn[18]
  PIN fn[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 596.000 548.240 600.000 ;
    END
  END fn[19]
  PIN fn[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 596.000 44.240 600.000 ;
    END
  END fn[1]
  PIN fn[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 596.000 576.240 600.000 ;
    END
  END fn[20]
  PIN fn[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 603.680 596.000 604.240 600.000 ;
    END
  END fn[21]
  PIN fn[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 596.000 632.240 600.000 ;
    END
  END fn[22]
  PIN fn[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 596.000 660.240 600.000 ;
    END
  END fn[23]
  PIN fn[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 596.000 688.240 600.000 ;
    END
  END fn[24]
  PIN fn[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 596.000 716.240 600.000 ;
    END
  END fn[25]
  PIN fn[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 596.000 744.240 600.000 ;
    END
  END fn[26]
  PIN fn[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 596.000 772.240 600.000 ;
    END
  END fn[27]
  PIN fn[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 596.000 800.240 600.000 ;
    END
  END fn[28]
  PIN fn[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 827.680 596.000 828.240 600.000 ;
    END
  END fn[29]
  PIN fn[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 596.000 72.240 600.000 ;
    END
  END fn[2]
  PIN fn[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 855.680 596.000 856.240 600.000 ;
    END
  END fn[30]
  PIN fn[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 596.000 884.240 600.000 ;
    END
  END fn[31]
  PIN fn[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 596.000 100.240 600.000 ;
    END
  END fn[3]
  PIN fn[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 596.000 128.240 600.000 ;
    END
  END fn[4]
  PIN fn[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 596.000 156.240 600.000 ;
    END
  END fn[5]
  PIN fn[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 596.000 184.240 600.000 ;
    END
  END fn[6]
  PIN fn[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 596.000 212.240 600.000 ;
    END
  END fn[7]
  PIN fn[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 596.000 240.240 600.000 ;
    END
  END fn[8]
  PIN fn[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 596.000 268.240 600.000 ;
    END
  END fn[9]
  PIN n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.480 0.000 47.040 4.000 ;
    END
  END n[0]
  PIN n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.080 0.000 136.640 4.000 ;
    END
  END n[1]
  PIN n[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.680 0.000 226.240 4.000 ;
    END
  END n[2]
  PIN n[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.280 0.000 315.840 4.000 ;
    END
  END n[3]
  PIN n[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 404.880 0.000 405.440 4.000 ;
    END
  END n[4]
  PIN n[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 494.480 0.000 495.040 4.000 ;
    END
  END n[5]
  PIN n[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.080 0.000 584.640 4.000 ;
    END
  END n[6]
  PIN n[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 673.680 0.000 674.240 4.000 ;
    END
  END n[7]
  PIN st
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 852.880 0.000 853.440 4.000 ;
    END
  END st
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 584.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 893.200 585.050 ;
      LAYER Metal2 ;
        RECT 16.540 595.700 43.380 596.000 ;
        RECT 44.540 595.700 71.380 596.000 ;
        RECT 72.540 595.700 99.380 596.000 ;
        RECT 100.540 595.700 127.380 596.000 ;
        RECT 128.540 595.700 155.380 596.000 ;
        RECT 156.540 595.700 183.380 596.000 ;
        RECT 184.540 595.700 211.380 596.000 ;
        RECT 212.540 595.700 239.380 596.000 ;
        RECT 240.540 595.700 267.380 596.000 ;
        RECT 268.540 595.700 295.380 596.000 ;
        RECT 296.540 595.700 323.380 596.000 ;
        RECT 324.540 595.700 351.380 596.000 ;
        RECT 352.540 595.700 379.380 596.000 ;
        RECT 380.540 595.700 407.380 596.000 ;
        RECT 408.540 595.700 435.380 596.000 ;
        RECT 436.540 595.700 463.380 596.000 ;
        RECT 464.540 595.700 491.380 596.000 ;
        RECT 492.540 595.700 519.380 596.000 ;
        RECT 520.540 595.700 547.380 596.000 ;
        RECT 548.540 595.700 575.380 596.000 ;
        RECT 576.540 595.700 603.380 596.000 ;
        RECT 604.540 595.700 631.380 596.000 ;
        RECT 632.540 595.700 659.380 596.000 ;
        RECT 660.540 595.700 687.380 596.000 ;
        RECT 688.540 595.700 715.380 596.000 ;
        RECT 716.540 595.700 743.380 596.000 ;
        RECT 744.540 595.700 771.380 596.000 ;
        RECT 772.540 595.700 799.380 596.000 ;
        RECT 800.540 595.700 827.380 596.000 ;
        RECT 828.540 595.700 855.380 596.000 ;
        RECT 856.540 595.700 883.380 596.000 ;
        RECT 884.540 595.700 884.660 596.000 ;
        RECT 15.820 4.300 884.660 595.700 ;
        RECT 15.820 4.000 46.180 4.300 ;
        RECT 47.340 4.000 135.780 4.300 ;
        RECT 136.940 4.000 225.380 4.300 ;
        RECT 226.540 4.000 314.980 4.300 ;
        RECT 316.140 4.000 404.580 4.300 ;
        RECT 405.740 4.000 494.180 4.300 ;
        RECT 495.340 4.000 583.780 4.300 ;
        RECT 584.940 4.000 673.380 4.300 ;
        RECT 674.540 4.000 762.980 4.300 ;
        RECT 764.140 4.000 852.580 4.300 ;
        RECT 853.740 4.000 884.660 4.300 ;
      LAYER Metal3 ;
        RECT 22.330 14.140 881.350 585.060 ;
      LAYER Metal4 ;
        RECT 369.740 41.530 405.940 563.270 ;
        RECT 408.140 41.530 408.660 563.270 ;
  END
END fibonacci
END LIBRARY

