* NGSPICE file created from fibonacci.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

.subckt fibonacci clk fn[0] fn[10] fn[11] fn[12] fn[13] fn[14] fn[15] fn[16] fn[17]
+ fn[18] fn[19] fn[1] fn[20] fn[21] fn[22] fn[23] fn[24] fn[25] fn[26] fn[27] fn[28]
+ fn[29] fn[2] fn[30] fn[31] fn[3] fn[4] fn[5] fn[6] fn[7] fn[8] fn[9] n[0] n[1] n[2]
+ n[3] n[4] n[5] n[6] n[7] st vdd vss
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_501_ _152_ _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_432_ c\[2\] c\[3\] _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__722__A1 _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_964_ _090_ net1 b\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_895_ _031_ net1 a\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_680_ _265_ _267_ _245_ _268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__437__I presente\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_947_ _073_ net1 b\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_878_ _014_ net1 a\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__447__A3 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_801_ _218_ _172_ _373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__438__A3 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__867__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_732_ _311_ _305_ _312_ _313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_663_ _250_ _252_ _253_ _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_594_ a\[15\] net17 _202_ _206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput31 net31 fn[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput20 net20 fn[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput42 net42 fn[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_715_ _275_ _294_ _298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_646_ a\[2\] b\[2\] _239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_577_ _196_ _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__561__S _187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_500_ b\[7\] _151_ _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__905__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_431_ c\[0\] _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_629_ _227_ _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__928__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__789__A2 _357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_963_ _089_ net1 b\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_894_ _030_ net1 a\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__689__A1 _274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_946_ _072_ net1 b\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_877_ _013_ net1 a\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__852__A1 _360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__538__I _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_800_ a\[23\] b\[23\] _372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_731_ a\[13\] b\[13\] _312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_662_ _250_ _252_ _245_ _253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_593_ _205_ _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_929_ _055_ net1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__961__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__825__A1 a\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput32 net32 fn[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput21 net21 fn[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__816__A1 a\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_714_ a\[11\] b\[11\] _286_ _294_ _296_ _297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_645_ _232_ _233_ _237_ _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_576_ a\[7\] net40 _192_ _196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__641__I _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I n[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__594__I0 a\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_430_ _098_ _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_628_ a\[28\] net31 _226_ _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_559_ _185_ _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__567__S _187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_962_ _088_ net1 b\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_893_ _029_ net1 a\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__918__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__689__A2 _275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_945_ _071_ net1 b\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_876_ _012_ net1 a\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__890__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_730_ a\[12\] b\[12\] _311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_661_ _251_ _252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_592_ a\[14\] net16 _202_ _205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_928_ _054_ net1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_859_ _418_ _422_ _423_ _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput33 net33 fn[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput22 net22 fn[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput11 net11 fn[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_713_ _295_ _296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_644_ a\[1\] b\[1\] _237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_575_ _195_ _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__951__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_627_ _208_ _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_558_ presente\[1\] _096_ _185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_489_ _124_ _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__567__I1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__716__A1 _280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__583__S _197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_961_ _087_ net1 b\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_892_ _028_ net1 a\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__630__I0 a\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_944_ _070_ net1 b\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_875_ _011_ net1 a\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__621__I0 a\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__908__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_660_ a\[4\] b\[4\] _251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_591_ _204_ _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__531__A2 _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_927_ _053_ net1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_858_ _418_ _422_ _124_ _423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_789_ _347_ _357_ _362_ _363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__513__A2 _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput34 net34 fn[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput23 net23 fn[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput12 net12 fn[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_712_ a\[11\] b\[11\] a\[10\] b\[10\] _295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_643_ _232_ _233_ _236_ _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__880__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_574_ a\[6\] net39 _192_ _195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__504__A2 _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__440__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_626_ _225_ _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_557_ _184_ _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_488_ _144_ _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_609_ a\[20\] net23 _215_ _216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__941__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_960_ _086_ net1 b\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_891_ _027_ net1 a\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__964__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__594__S _202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__630__I1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__846__A1 _411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_943_ _069_ net1 b\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_874_ _010_ net1 a\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_590_ a\[13\] net15 _202_ _204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_926_ _052_ net1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_857_ _415_ _419_ _420_ _411_ _421_ _422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_788_ a\[20\] b\[20\] _362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 net24 fn[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput13 net13 fn[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput35 net35 fn[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_711_ _284_ _291_ _294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_642_ _232_ _233_ _235_ _236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_573_ _194_ _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_909_ _035_ net1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__440__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__579__I0 a\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_625_ a\[27\] net30 _221_ _225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_556_ b\[31\] _099_ _184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_487_ b\[2\] _141_ _144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__870__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_608_ _208_ _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_539_ b\[23\] _174_ _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__893__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_890_ _026_ net1 a\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__791__A1 _360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_942_ _068_ net1 b\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_873_ _009_ net1 a\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__782__A1 _330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__931__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__954__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_925_ _051_ net1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__489__I _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_856_ a\[29\] b\[29\] _421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_787_ a\[21\] b\[21\] _361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__746__A1 a\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput25 net25 fn[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput14 net14 fn[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_135_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput36 net36 fn[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_710_ _290_ _291_ _293_ _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_641_ _234_ _235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_572_ a\[5\] net38 _192_ _194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_908_ _034_ net1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_839_ a\[24\] b\[24\] _387_ _406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__440__A3 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_624_ _224_ _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_555_ _183_ _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_486_ _143_ _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__587__I _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_607_ _214_ _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_538_ _098_ _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_469_ c\[4\] _126_ _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__552__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__814__B _358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__543__A2 _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_941_ _067_ net1 b\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_872_ _008_ net1 a\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__883__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__782__A2 _350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__461__A1 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_924_ _050_ net1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_855_ _412_ _414_ _420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_786_ _133_ _360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__452__A1 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput15 net15 fn[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput26 net26 fn[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput37 net37 fn[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_640_ _097_ _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_571_ _193_ _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__921__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__673__A1 a\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_907_ _033_ net1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_838_ _401_ _404_ _405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_769_ a\[19\] b\[19\] _345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__440__A4 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__944__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_623_ a\[26\] net29 _221_ _224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__783__I _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_554_ b\[30\] _179_ _183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_485_ b\[1\] _141_ _143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__967__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__642__B _235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__637__A1 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_606_ a\[19\] net21 _209_ _214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__727__B _292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_537_ _173_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_468_ _114_ _129_ _130_ c1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__598__I _208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_940_ _066_ net1 b\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_871_ _007_ net1 a\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_923_ _049_ net1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_854_ a\[29\] b\[29\] _419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__786__I _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_785_ _347_ _357_ _359_ _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__873__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput27 net27 fn[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput16 net16 fn[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput38 net38 fn[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_570_ a\[4\] net37 _192_ _193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_906_ _032_ net1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_837_ _384_ _386_ _388_ _394_ _404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_768_ _338_ _341_ _343_ _344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_699_ a\[10\] b\[10\] _284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__896__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_622_ _223_ _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_553_ _182_ _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_484_ _142_ _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__911__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_605_ _213_ _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__800__A2 b\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_536_ _172_ _168_ _173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_467_ net6 _117_ _130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__934__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__957__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_519_ _162_ _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_870_ _006_ net1 a\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__749__A1 _297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_922_ _048_ net1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_853_ a\[30\] b\[30\] _418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_784_ _347_ _357_ _358_ _359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 fn[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput17 net17 fn[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput39 net39 fn[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_905_ c1\[7\] net1 c\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_836_ _283_ _402_ _403_ _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_767_ a\[18\] b\[18\] _343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_698_ _113_ _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__611__S _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_621_ a\[25\] net28 _221_ _223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_552_ b\[29\] _179_ _182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_483_ b\[0\] _141_ _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_819_ _386_ _388_ _389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__476__B _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__606__S _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__886__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_604_ a\[18\] net20 _209_ _213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_535_ b\[22\] _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_466_ c\[4\] _126_ _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__785__A2 _357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_518_ b\[15\] _161_ _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__901__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_449_ _113_ _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__464__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__924__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__947__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__614__S _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_921_ _047_ net1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_852_ _360_ _417_ _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_783_ _234_ _358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__428__A1 presente\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput29 net29 fn[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput18 net18 fn[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__667__A1 a\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__609__S _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_904_ c1\[6\] net1 c\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_835_ _400_ _398_ _401_ _403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__830__A1 _235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_766_ _338_ _341_ _342_ _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_697_ _254_ _282_ _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__821__A1 _383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_620_ _222_ _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__812__A1 _329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_551_ _181_ _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_482_ _098_ _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_818_ _387_ _388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_749_ _297_ _323_ _325_ _326_ _327_ _328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_603_ _212_ _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_534_ _171_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_465_ _128_ c1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__572__I0 a\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_517_ _150_ _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_448_ _114_ _105_ _115_ _110_ futuro\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__876__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__680__B _245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__464__A2 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__765__B _292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__899__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__675__B _245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__630__S _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_920_ _046_ net1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_851_ _414_ _416_ _417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_782_ _330_ _350_ _356_ _357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__428__A2 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 net19 fn[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__914__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_903_ c1\[5\] net1 c\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_834_ _400_ _398_ _401_ _402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_765_ _338_ _341_ _292_ _342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_696_ _280_ _281_ _282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_1_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__937__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__812__A2 _350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_550_ b\[28\] _179_ _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_481_ _114_ _139_ _140_ c1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_817_ a\[25\] b\[25\] _387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_748_ _313_ _322_ _327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_679_ a\[6\] b\[6\] _266_ _267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__558__A1 presente\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__858__B _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_602_ _211_ net19 _209_ _212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__797__A1 _357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_533_ b\[21\] _168_ _171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_464_ net5 _099_ _127_ _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__563__I1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_516_ _160_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_447_ net10 _106_ _096_ _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__517__I _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__628__S _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_850_ _411_ _412_ _415_ _416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_781_ _352_ _355_ _356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__866__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__889__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_902_ c1\[4\] net1 c\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_833_ a\[27\] b\[27\] _401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_764_ _211_ _165_ _334_ _340_ _341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_695_ a\[8\] b\[8\] _276_ _281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input8_I n[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_480_ net9 _133_ _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__500__A2 _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_816_ a\[25\] b\[25\] _386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_747_ a\[15\] b\[15\] _326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_678_ _258_ _263_ _266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__904__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__558__A2 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__927__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_601_ a\[17\] _211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__797__A2 _366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_532_ _170_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_463_ _124_ _125_ _126_ _127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__784__B _358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_515_ b\[14\] _156_ _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_446_ _113_ _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__458__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__697__A1 _254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__708__I _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__688__A1 a\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__860__A1 a\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__618__I _208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_429_ _097_ _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__679__A1 a\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 clk net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__528__I _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_780_ _343_ _353_ _354_ _355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__842__A1 a\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__833__A1 a\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__960__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_901_ c1\[3\] net1 c\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_832_ a\[26\] b\[26\] _400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__815__A1 _383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_763_ _339_ _340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_694_ _278_ _279_ _280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_815_ _383_ _384_ _385_ _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_746_ a\[15\] b\[15\] _317_ _325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_677_ a\[7\] b\[7\] _265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__879__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__494__A2 _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_600_ _210_ _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_531_ b\[20\] _168_ _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_462_ c\[0\] c\[1\] _101_ _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_144_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__446__I _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__485__A2 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_729_ a\[14\] b\[14\] _310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__467__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_514_ _159_ _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_445_ _112_ _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__458__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__917__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_428_ presente\[1\] _096_ _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 n[0] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__565__S _187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_900_ c1\[2\] net1 c\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_831_ _395_ _397_ _399_ _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_762_ a\[16\] b\[16\] a\[17\] b\[17\] _339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__449__I _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_693_ a\[9\] b\[9\] _279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__806__A2 _366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_814_ _383_ _384_ _358_ _385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_745_ _280_ _298_ _323_ _324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_676_ _258_ _263_ _264_ _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__950__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__715__A1 _275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_530_ _169_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_461_ _100_ _103_ c\[2\] c\[3\] _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__706__A1 a\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_728_ _307_ _308_ _309_ _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_659_ a\[3\] b\[3\] _238_ _247_ _249_ _250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__547__I _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_513_ b\[13\] _156_ _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_444_ _106_ presente\[0\] _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__869__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_427_ presente\[0\] _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 n[1] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__560__I _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__907__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__581__S _197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__521__A2 _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_830_ _235_ _398_ _399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_761_ _337_ _338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_692_ a\[9\] b\[9\] _278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_959_ _085_ net1 b\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_813_ a\[24\] b\[24\] _384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_744_ _302_ _305_ _306_ _322_ _323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_675_ _258_ _263_ _245_ _264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I n[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__651__A1 _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_460_ _097_ _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_727_ _307_ _308_ _292_ _309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_658_ _242_ _248_ _249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_589_ _203_ _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__653__I _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_512_ _158_ _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__940__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_443_ _111_ futuro\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__863__A1 _360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__854__A1 a\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__963__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__579__S _197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__836__A1 _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 n[2] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__827__A1 a\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__751__I _329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__700__B a\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_760_ a\[18\] b\[18\] _337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_691_ _276_ _277_ _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_958_ _084_ net1 b\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_889_ _025_ net1 a\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__592__S _202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_812_ _329_ _350_ _377_ _381_ _382_ _383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_743_ _310_ _318_ _322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_674_ _255_ _261_ _262_ _263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_726_ a\[12\] b\[12\] _304_ _308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_657_ a\[3\] b\[3\] _248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_588_ a\[12\] net14 _202_ _203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__892__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_511_ b\[12\] _156_ _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_442_ _099_ _105_ _107_ _110_ _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_709_ _290_ _291_ _292_ _293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__664__I _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__781__A1 _352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput5 n[3] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__930__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__569__I _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__754__A1 _330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__953__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__809__A2 _379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__745__A1 _280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_690_ _274_ _275_ _235_ _277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__736__A1 _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_957_ _083_ net1 b\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_888_ _024_ net1 a\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__718__A1 _297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_811_ a\[23\] b\[23\] _382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_742_ _321_ _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_673_ a\[5\] b\[5\] _262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_725_ _305_ _306_ _307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_656_ _239_ _241_ _247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_587_ _186_ _202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_510_ _157_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__632__I0 a\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_441_ _108_ _109_ _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_708_ _234_ _292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__623__I0 a\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_639_ a\[1\] b\[1\] _233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__804__B _358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__533__A2 _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 n[4] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__882__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__524__A2 _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__515__A2 _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__709__B _292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__451__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__506__A2 _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__690__A1 _274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__442__A1 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_956_ _082_ net1 b\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_887_ _023_ net1 a\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__920__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__663__A1 _250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_810_ _218_ _172_ a\[23\] b\[23\] _380_ _381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_741_ _099_ _319_ _320_ _321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_672_ _259_ _260_ _261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__943__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_939_ _065_ net1 b\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__966__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_724_ a\[13\] b\[13\] _306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_655_ _241_ _244_ _246_ _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_586_ _201_ _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I n[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__857__B2 _411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__632__I1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_440_ net9 net8 net2 net3 _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__848__A1 a\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_707_ a\[11\] b\[11\] _291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_638_ a\[0\] b\[0\] _232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_569_ _186_ _192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 n[5] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__451__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__690__A2 _275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__872__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_955_ _081_ net1 b\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_886_ _022_ net1 a\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput10 st net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__895__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_740_ _317_ _316_ _318_ _320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_671_ a\[5\] b\[5\] _260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_938_ _064_ net1 b\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_869_ _005_ net1 a\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__823__B _358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__910__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_723_ a\[13\] b\[13\] _305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_654_ _241_ _244_ _245_ _246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_585_ a\[11\] net13 _197_ _201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__933__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_706_ a\[10\] b\[10\] _289_ _290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_637_ _141_ _231_ _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_568_ _191_ _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_499_ _150_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__536__A1 _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__956__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput8 n[6] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_954_ _080_ net1 b\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_885_ _021_ net1 a\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_670_ a\[4\] b\[4\] _259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_937_ _063_ net1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_868_ _004_ net1 a\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_799_ _360_ _371_ _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_722_ _283_ _303_ _304_ _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_653_ _234_ _245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_584_ _200_ _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__885__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__554__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__545__A2 _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_705_ _283_ _288_ _289_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_636_ a\[0\] b\[0\] _231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_567_ a\[3\] net36 _187_ _191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__784__A2 _357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__536__A2 _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_498_ _097_ _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__472__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__654__B _245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__900__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__463__A1 _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__518__A2 _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__454__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 n[7] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_619_ a\[24\] net27 _221_ _222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__923__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__509__A2 _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__604__S _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__684__A1 a\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__946__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__436__A1 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__969__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_953_ _079_ net1 b\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_884_ _020_ net1 a\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__648__A1 _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__662__B _245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output11_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_936_ _062_ net1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_867_ _003_ net1 a\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_798_ _365_ _370_ _371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_721_ _301_ _302_ _304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_652_ _242_ _243_ _244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_583_ a\[10\] net12 _197_ _200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_919_ _045_ net1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__490__A2 _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I st vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_704_ _284_ _287_ _289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_635_ _230_ _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_566_ _190_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_497_ _149_ _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I n[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__472__A2 _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__875__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__454__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_618_ _208_ _221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_549_ _180_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__898__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__913__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_952_ _078_ net1 b\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_883_ _019_ net1 a\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__936__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__811__A2 b\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_935_ _061_ net1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_866_ _002_ net1 a\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__802__A2 _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_797_ _357_ _366_ _369_ _370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__959__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_720_ _301_ _302_ _303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_651_ _238_ _239_ _243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_582_ _199_ _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_918_ _044_ net1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_849_ a\[28\] b\[28\] _415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__539__A1 b\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_703_ _284_ _287_ _288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_634_ a\[31\] net35 _226_ _230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_565_ a\[2\] net33 _187_ _190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_496_ b\[6\] _145_ _149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__463__A3 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_617_ _220_ _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_548_ b\[27\] _179_ _180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_479_ c\[7\] _138_ _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__865__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__430__I _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_951_ _077_ net1 b\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_882_ _018_ net1 a\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__888__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_934_ _060_ net1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_865_ _001_ net1 a\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_796_ _367_ _368_ _369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__903__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_650_ a\[2\] b\[2\] _242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_581_ a\[9\] net42 _197_ _199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__548__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_917_ _043_ net1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_848_ a\[29\] b\[29\] _414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__926__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_779_ a\[19\] b\[19\] _354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__539__A2 _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__949__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_702_ _276_ _279_ _286_ _287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_633_ _229_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_564_ _189_ _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_495_ _148_ _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__696__A1 _280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__634__S _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__687__A1 _250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__439__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_616_ a\[23\] net26 _215_ _220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__608__I _208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_547_ _098_ _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_478_ _102_ _121_ _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__850__A1 _411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__669__A1 a\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__841__A1 a\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__832__A1 a\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_950_ _076_ net1 b\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_881_ _017_ net1 a\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__814__A1 _383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__583__I0 a\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_933_ _059_ net1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_864_ _000_ net1 a\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_795_ a\[21\] b\[21\] a\[20\] b\[20\] _368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__574__I0 a\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_580_ _198_ _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__878__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_916_ _042_ net1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_847_ _411_ _412_ _413_ _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_778_ a\[19\] b\[19\] _353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__466__A2 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_701_ _278_ _285_ _286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_632_ a\[30\] net34 _226_ _229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_563_ a\[1\] net22 _187_ _189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_494_ b\[5\] _145_ _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__916__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__439__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_615_ _219_ _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_546_ _178_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_477_ _135_ _116_ _136_ _137_ c1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__939__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_529_ b\[19\] _168_ _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_880_ _016_ net1 a\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__750__A1 _274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__741__A1 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_932_ _058_ net1 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_863_ _360_ _426_ _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__799__A1 _360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_794_ a\[21\] b\[21\] _367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__565__I1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__705__A1 _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_915_ _041_ net1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_846_ _411_ _412_ _124_ _413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_777_ _351_ _337_ _339_ _345_ _352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__627__I _208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__563__S _187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__475__A3 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_700_ a\[9\] b\[9\] a\[8\] b\[8\] _285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_631_ _228_ _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_562_ _188_ _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_493_ _147_ _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_829_ _396_ _392_ _394_ _388_ _398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__868__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_614_ _218_ net25 _215_ _219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_545_ b\[26\] _174_ _178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_476_ _102_ _121_ _113_ _137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_528_ _150_ _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_459_ _116_ _122_ _123_ c1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__906__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__511__A2 _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__502__A2 _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__929__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_931_ _057_ net1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_862_ a\[31\] b\[31\] _425_ _426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_793_ _347_ _361_ _366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_914_ _040_ net1 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_845_ a\[28\] b\[28\] _412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_134_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_776_ _211_ _165_ _351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__699__A1 a\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_630_ a\[29\] net32 _226_ _228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_561_ a\[0\] net11 _187_ _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_492_ b\[4\] _145_ _147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__862__A1 a\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_828_ _396_ _392_ _388_ _397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_759_ _254_ _336_ _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__853__A1 a\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__439__A4 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__844__A1 _383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__962__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_613_ a\[22\] _218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_544_ _177_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_475_ c\[4\] c\[5\] _126_ c\[6\] _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__817__A1 a\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_527_ _167_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_458_ net4 _117_ _123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__808__A1 _352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_930_ _056_ net1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__496__A2 _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_861_ _418_ _422_ _424_ _425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_792_ a\[22\] b\[22\] _365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__487__A2 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__919__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__469__A2 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_913_ _039_ net1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_844_ _383_ _405_ _407_ _410_ _411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_134_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_775_ _348_ _333_ _349_ _350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_560_ _186_ _187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_491_ _146_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__891__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_827_ a\[25\] b\[25\] _396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_758_ _333_ _335_ _336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_689_ _274_ _275_ _276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__590__S _202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_612_ _217_ _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_543_ b\[25\] _174_ _177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_474_ net8 _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__474__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__585__S _197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__771__A1 _254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_526_ b\[18\] _161_ _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_457_ c\[2\] _121_ _122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__753__A1 _330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__952__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_509_ b\[11\] _156_ _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__717__A1 _274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_860_ a\[30\] b\[30\] _424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_791_ _360_ _364_ _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__482__I _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_912_ _038_ net1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_843_ _400_ _408_ _409_ _410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_774_ _338_ _345_ _349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__588__S _202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I n[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_490_ b\[3\] _145_ _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_826_ _394_ _395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_757_ _207_ _163_ _334_ _335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_688_ a\[8\] b\[8\] _275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__550__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__909__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__541__A2 _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_611_ a\[21\] net24 _215_ _217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_542_ _176_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_473_ _114_ _132_ _134_ c1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_809_ _378_ _379_ _373_ _380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__881__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_525_ _166_ _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_456_ c\[0\] _103_ _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__671__A1 a\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_508_ _150_ _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_439_ net4 net5 net6 net7 _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__662__A1 _250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_790_ _361_ _363_ _364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__712__B a\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__942__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_911_ _037_ net1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_842_ a\[27\] b\[27\] _409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__965__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_773_ _207_ _163_ _348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__856__A1 a\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__578__I _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__847__A1 _411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_825_ a\[26\] b\[26\] _394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_756_ _330_ _331_ _334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_687_ _250_ _270_ _271_ _272_ _273_ _274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__599__S _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_610_ _216_ _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_541_ b\[24\] _174_ _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_472_ net7 _133_ _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_808_ _352_ _355_ _366_ _379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_739_ _317_ _316_ _318_ _319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_524_ _165_ _161_ _166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_455_ _116_ _119_ _120_ c1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_507_ _155_ _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_438_ net10 _106_ _096_ _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__871__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__894__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_910_ _036_ net1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_841_ a\[27\] b\[27\] _408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_772_ a\[20\] b\[20\] _347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__808__B _366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__932__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_824_ _389_ _392_ _393_ _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_755_ _211_ _165_ _333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_686_ _262_ _261_ _269_ _273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__955__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_540_ _175_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_471_ _112_ _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__499__I _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_807_ _369_ _378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_738_ a\[15\] b\[15\] _318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_669_ a\[6\] b\[6\] _258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__756__A1 _330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__747__A1 a\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_523_ b\[17\] _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__738__A1 a\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_454_ net3 _117_ _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_506_ b\[10\] _151_ _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_437_ presente\[1\] _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_840_ _386_ _406_ _401_ _395_ _407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_134_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_771_ _254_ _346_ _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__634__I0 a\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_969_ _095_ net1 b\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__625__I0 a\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__884__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_823_ _389_ _392_ _358_ _393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_754_ _330_ _331_ _332_ _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__480__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_685_ a\[7\] b\[7\] _272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I n[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__526__A2 _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_470_ c\[5\] _131_ _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_806_ _365_ _366_ _372_ _377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__453__A1 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_737_ a\[14\] b\[14\] _317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_668_ _254_ _257_ _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_599_ _207_ net18 _209_ _210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__922__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_522_ _164_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_453_ _100_ _103_ _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__945__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__665__A1 _250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__968__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_505_ _154_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_436_ _100_ _102_ _104_ _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__647__A1 _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__810__B2 b\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__698__I _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__647__B _235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__602__S _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_770_ _344_ _345_ _346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__634__I1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_968_ _094_ net1 b\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_899_ c1\[1\] net1 c\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__625__I1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__616__I1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_822_ _390_ _391_ _392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_753_ _330_ _331_ _292_ _332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__480__A2 _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_684_ a\[6\] b\[6\] a\[7\] b\[7\] _271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_805_ _372_ _375_ _376_ _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_736_ _283_ _314_ _316_ _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_667_ a\[5\] b\[5\] _256_ _257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_598_ _208_ _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__874__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_521_ _163_ _161_ _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_452_ _100_ _116_ _118_ c1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__897__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_719_ a\[12\] b\[12\] _302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_504_ b\[9\] _151_ _154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_435_ _103_ c\[7\] _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__912__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__810__A2 _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__935__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__801__A2 _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__753__B _292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__958__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__570__I1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_967_ _093_ net1 b\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_898_ c1\[0\] net1 c\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__561__I1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_821_ _383_ _384_ _391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_752_ _207_ _163_ _331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_683_ _251_ _260_ _262_ _269_ _270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__759__A1 _254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_804_ _372_ _375_ _358_ _376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_735_ _305_ _308_ _315_ _312_ _316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_666_ a\[4\] b\[4\] _255_ _256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_597_ _185_ _208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_520_ b\[16\] _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__846__B _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_451_ net2 _117_ _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__659__B1 _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_718_ _297_ _300_ _301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_649_ a\[3\] b\[3\] _241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__864__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_503_ _153_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_434_ c\[1\] _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__887__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__616__S _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__556__A2 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__902__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_966_ _092_ net1 b\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_897_ futuro\[1\] net1 presente\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__925__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__529__A2 _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_820_ a\[24\] b\[24\] _390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_751_ _329_ _330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_682_ _258_ _265_ _269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__948__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_949_ _075_ net1 b\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__695__A1 a\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__447__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__438__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_803_ _373_ _370_ _374_ _375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_734_ _310_ _315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_665_ _250_ _252_ _255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_596_ a\[16\] _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I n[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__508__I _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__668__A1 _254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_450_ _112_ _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput40 net40 fn[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_717_ _274_ _299_ _300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_648_ _238_ _239_ _240_ _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_579_ a\[8\] net41 _197_ _198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_502_ b\[8\] _151_ _153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_433_ c\[4\] c\[5\] c\[6\] _101_ _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__632__S _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__492__A2 _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__483__A2 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_965_ _091_ net1 b\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_896_ futuro\[0\] net1 presente\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__877__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__690__B _235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_750_ _274_ _324_ _328_ _329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_681_ _265_ _267_ _268_ _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_948_ _074_ net1 b\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_879_ _015_ net1 a\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_802_ _218_ _172_ _374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_733_ _304_ _306_ _310_ _313_ _314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_664_ _133_ _254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_595_ _206_ _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__915__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__938__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput30 net30 fn[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput41 net41 fn[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_716_ _280_ _298_ _299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_647_ _238_ _239_ _235_ _240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_578_ _186_ _197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

