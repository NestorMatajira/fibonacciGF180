magic
tech gf180mcuC
magscale 1 10
timestamp 1670116059
<< metal1 >>
rect 158162 117070 158174 117122
rect 158226 117119 158238 117122
rect 159282 117119 159294 117122
rect 158226 117073 159294 117119
rect 158226 117070 158238 117073
rect 159282 117070 159294 117073
rect 159346 117070 159358 117122
rect 30482 116958 30494 117010
rect 30546 117007 30558 117010
rect 31602 117007 31614 117010
rect 30546 116961 31614 117007
rect 30546 116958 30558 116961
rect 31602 116958 31614 116961
rect 31666 116958 31678 117010
rect 77522 116958 77534 117010
rect 77586 117007 77598 117010
rect 78642 117007 78654 117010
rect 77586 116961 78654 117007
rect 77586 116958 77598 116961
rect 78642 116958 78654 116961
rect 78706 116958 78718 117010
rect 111122 116958 111134 117010
rect 111186 117007 111198 117010
rect 112242 117007 112254 117010
rect 111186 116961 112254 117007
rect 111186 116958 111198 116961
rect 112242 116958 112254 116961
rect 112306 116958 112318 117010
rect 112690 116958 112702 117010
rect 112754 117007 112766 117010
rect 113586 117007 113598 117010
rect 112754 116961 113598 117007
rect 112754 116958 112766 116961
rect 113586 116958 113598 116961
rect 113650 116958 113662 117010
rect 134642 116958 134654 117010
rect 134706 117007 134718 117010
rect 135762 117007 135774 117010
rect 134706 116961 135774 117007
rect 134706 116958 134718 116961
rect 135762 116958 135774 116961
rect 135826 116958 135838 117010
rect 136210 116958 136222 117010
rect 136274 117007 136286 117010
rect 137554 117007 137566 117010
rect 136274 116961 137566 117007
rect 136274 116958 136286 116961
rect 137554 116958 137566 116961
rect 137618 116958 137630 117010
rect 159730 116958 159742 117010
rect 159794 117007 159806 117010
rect 160402 117007 160414 117010
rect 159794 116961 160414 117007
rect 159794 116958 159806 116961
rect 160402 116958 160414 116961
rect 160466 116958 160478 117010
rect 1344 116842 178640 116876
rect 1344 116790 4478 116842
rect 4530 116790 4582 116842
rect 4634 116790 4686 116842
rect 4738 116790 35198 116842
rect 35250 116790 35302 116842
rect 35354 116790 35406 116842
rect 35458 116790 65918 116842
rect 65970 116790 66022 116842
rect 66074 116790 66126 116842
rect 66178 116790 96638 116842
rect 96690 116790 96742 116842
rect 96794 116790 96846 116842
rect 96898 116790 127358 116842
rect 127410 116790 127462 116842
rect 127514 116790 127566 116842
rect 127618 116790 158078 116842
rect 158130 116790 158182 116842
rect 158234 116790 158286 116842
rect 158338 116790 178640 116842
rect 1344 116756 178640 116790
rect 3378 116510 3390 116562
rect 3442 116510 3454 116562
rect 5954 116510 5966 116562
rect 6018 116510 6030 116562
rect 8418 116510 8430 116562
rect 8482 116510 8494 116562
rect 10098 116510 10110 116562
rect 10162 116510 10174 116562
rect 14354 116510 14366 116562
rect 14418 116510 14430 116562
rect 19058 116510 19070 116562
rect 19122 116510 19134 116562
rect 22194 116510 22206 116562
rect 22258 116510 22270 116562
rect 23538 116510 23550 116562
rect 23602 116510 23614 116562
rect 27346 116510 27358 116562
rect 27410 116510 27422 116562
rect 29474 116510 29486 116562
rect 29538 116510 29550 116562
rect 31938 116510 31950 116562
rect 32002 116510 32014 116562
rect 33618 116510 33630 116562
rect 33682 116510 33694 116562
rect 37874 116510 37886 116562
rect 37938 116510 37950 116562
rect 42578 116510 42590 116562
rect 42642 116510 42654 116562
rect 45714 116510 45726 116562
rect 45778 116510 45790 116562
rect 47058 116510 47070 116562
rect 47122 116510 47134 116562
rect 50866 116510 50878 116562
rect 50930 116510 50942 116562
rect 52994 116510 53006 116562
rect 53058 116510 53070 116562
rect 55458 116510 55470 116562
rect 55522 116510 55534 116562
rect 57138 116510 57150 116562
rect 57202 116510 57214 116562
rect 61394 116510 61406 116562
rect 61458 116510 61470 116562
rect 66098 116510 66110 116562
rect 66162 116510 66174 116562
rect 69234 116510 69246 116562
rect 69298 116510 69310 116562
rect 70578 116510 70590 116562
rect 70642 116510 70654 116562
rect 74386 116510 74398 116562
rect 74450 116510 74462 116562
rect 76514 116510 76526 116562
rect 76578 116510 76590 116562
rect 78978 116510 78990 116562
rect 79042 116510 79054 116562
rect 80658 116510 80670 116562
rect 80722 116510 80734 116562
rect 84914 116510 84926 116562
rect 84978 116510 84990 116562
rect 89618 116510 89630 116562
rect 89682 116510 89694 116562
rect 93202 116510 93214 116562
rect 93266 116510 93278 116562
rect 97906 116510 97918 116562
rect 97970 116510 97982 116562
rect 100034 116510 100046 116562
rect 100098 116510 100110 116562
rect 102498 116510 102510 116562
rect 102562 116510 102574 116562
rect 104178 116510 104190 116562
rect 104242 116510 104254 116562
rect 108322 116510 108334 116562
rect 108386 116510 108398 116562
rect 112242 116510 112254 116562
rect 112306 116510 112318 116562
rect 113586 116510 113598 116562
rect 113650 116510 113662 116562
rect 116722 116510 116734 116562
rect 116786 116510 116798 116562
rect 121426 116510 121438 116562
rect 121490 116510 121502 116562
rect 124002 116510 124014 116562
rect 124066 116510 124078 116562
rect 126018 116510 126030 116562
rect 126082 116510 126094 116562
rect 127922 116510 127934 116562
rect 127986 116510 127998 116562
rect 131842 116510 131854 116562
rect 131906 116510 131918 116562
rect 135762 116510 135774 116562
rect 135826 116510 135838 116562
rect 137554 116510 137566 116562
rect 137618 116510 137630 116562
rect 140242 116510 140254 116562
rect 140306 116510 140318 116562
rect 144946 116510 144958 116562
rect 145010 116510 145022 116562
rect 147522 116510 147534 116562
rect 147586 116510 147598 116562
rect 149538 116510 149550 116562
rect 149602 116510 149614 116562
rect 151442 116510 151454 116562
rect 151506 116510 151518 116562
rect 155362 116510 155374 116562
rect 155426 116510 155438 116562
rect 159282 116510 159294 116562
rect 159346 116510 159358 116562
rect 163762 116510 163774 116562
rect 163826 116510 163838 116562
rect 168466 116510 168478 116562
rect 168530 116510 168542 116562
rect 173058 116510 173070 116562
rect 173122 116510 173134 116562
rect 20526 116450 20578 116462
rect 81902 116450 81954 116462
rect 146078 116450 146130 116462
rect 4386 116398 4398 116450
rect 4450 116398 4462 116450
rect 6738 116398 6750 116450
rect 6802 116398 6814 116450
rect 7634 116398 7646 116450
rect 7698 116398 7710 116450
rect 10882 116398 10894 116450
rect 10946 116398 10958 116450
rect 15362 116398 15374 116450
rect 15426 116398 15438 116450
rect 19842 116398 19854 116450
rect 19906 116398 19918 116450
rect 21746 116398 21758 116450
rect 21810 116398 21822 116450
rect 24546 116398 24558 116450
rect 24610 116398 24622 116450
rect 26674 116398 26686 116450
rect 26738 116398 26750 116450
rect 30482 116398 30494 116450
rect 30546 116398 30558 116450
rect 31154 116398 31166 116450
rect 31218 116398 31230 116450
rect 34402 116398 34414 116450
rect 34466 116398 34478 116450
rect 38882 116398 38894 116450
rect 38946 116398 38958 116450
rect 43586 116398 43598 116450
rect 43650 116398 43662 116450
rect 45266 116398 45278 116450
rect 45330 116398 45342 116450
rect 48066 116398 48078 116450
rect 48130 116398 48142 116450
rect 50194 116398 50206 116450
rect 50258 116398 50270 116450
rect 53778 116398 53790 116450
rect 53842 116398 53854 116450
rect 54674 116398 54686 116450
rect 54738 116398 54750 116450
rect 57922 116398 57934 116450
rect 57986 116398 57998 116450
rect 62402 116398 62414 116450
rect 62466 116398 62478 116450
rect 67106 116398 67118 116450
rect 67170 116398 67182 116450
rect 68786 116398 68798 116450
rect 68850 116398 68862 116450
rect 71362 116398 71374 116450
rect 71426 116398 71438 116450
rect 73714 116398 73726 116450
rect 73778 116398 73790 116450
rect 77522 116398 77534 116450
rect 77586 116398 77598 116450
rect 78194 116398 78206 116450
rect 78258 116398 78270 116450
rect 81218 116398 81230 116450
rect 81282 116398 81294 116450
rect 85922 116398 85934 116450
rect 85986 116398 85998 116450
rect 90626 116398 90638 116450
rect 90690 116398 90702 116450
rect 92530 116398 92542 116450
rect 92594 116398 92606 116450
rect 97234 116398 97246 116450
rect 97298 116398 97310 116450
rect 101042 116398 101054 116450
rect 101106 116398 101118 116450
rect 101714 116398 101726 116450
rect 101778 116398 101790 116450
rect 104962 116398 104974 116450
rect 105026 116398 105038 116450
rect 107650 116398 107662 116450
rect 107714 116398 107726 116450
rect 111570 116398 111582 116450
rect 111634 116398 111646 116450
rect 114370 116398 114382 116450
rect 114434 116398 114446 116450
rect 116050 116398 116062 116450
rect 116114 116398 116126 116450
rect 120978 116398 120990 116450
rect 121042 116398 121054 116450
rect 123330 116398 123342 116450
rect 123394 116398 123406 116450
rect 125234 116398 125246 116450
rect 125298 116398 125310 116450
rect 127250 116398 127262 116450
rect 127314 116398 127326 116450
rect 131170 116398 131182 116450
rect 131234 116398 131246 116450
rect 135090 116398 135102 116450
rect 135154 116398 135166 116450
rect 136882 116398 136894 116450
rect 136946 116398 136958 116450
rect 139570 116398 139582 116450
rect 139634 116398 139646 116450
rect 144274 116398 144286 116450
rect 144338 116398 144350 116450
rect 146850 116398 146862 116450
rect 146914 116398 146926 116450
rect 148754 116398 148766 116450
rect 148818 116398 148830 116450
rect 150770 116398 150782 116450
rect 150834 116398 150846 116450
rect 154690 116398 154702 116450
rect 154754 116398 154766 116450
rect 158610 116398 158622 116450
rect 158674 116398 158686 116450
rect 163090 116398 163102 116450
rect 163154 116398 163166 116450
rect 167794 116398 167806 116450
rect 167858 116398 167870 116450
rect 172274 116398 172286 116450
rect 172338 116398 172350 116450
rect 20526 116386 20578 116398
rect 81902 116386 81954 116398
rect 146078 116386 146130 116398
rect 39342 116338 39394 116350
rect 39342 116274 39394 116286
rect 160414 116338 160466 116350
rect 160414 116274 160466 116286
rect 164894 116338 164946 116350
rect 164894 116274 164946 116286
rect 170382 116338 170434 116350
rect 170382 116274 170434 116286
rect 174302 116338 174354 116350
rect 174302 116274 174354 116286
rect 177214 116338 177266 116350
rect 177214 116274 177266 116286
rect 11342 116226 11394 116238
rect 11342 116162 11394 116174
rect 15822 116226 15874 116238
rect 15822 116162 15874 116174
rect 25230 116226 25282 116238
rect 25230 116162 25282 116174
rect 34862 116226 34914 116238
rect 34862 116162 34914 116174
rect 44046 116226 44098 116238
rect 44046 116162 44098 116174
rect 48750 116226 48802 116238
rect 48750 116162 48802 116174
rect 58382 116226 58434 116238
rect 58382 116162 58434 116174
rect 62862 116226 62914 116238
rect 62862 116162 62914 116174
rect 67566 116226 67618 116238
rect 67566 116162 67618 116174
rect 72270 116226 72322 116238
rect 72270 116162 72322 116174
rect 86382 116226 86434 116238
rect 86382 116162 86434 116174
rect 91086 116226 91138 116238
rect 91086 116162 91138 116174
rect 105422 116226 105474 116238
rect 105422 116162 105474 116174
rect 122558 116226 122610 116238
rect 122558 116162 122610 116174
rect 1344 116058 178640 116092
rect 1344 116006 19838 116058
rect 19890 116006 19942 116058
rect 19994 116006 20046 116058
rect 20098 116006 50558 116058
rect 50610 116006 50662 116058
rect 50714 116006 50766 116058
rect 50818 116006 81278 116058
rect 81330 116006 81382 116058
rect 81434 116006 81486 116058
rect 81538 116006 111998 116058
rect 112050 116006 112102 116058
rect 112154 116006 112206 116058
rect 112258 116006 142718 116058
rect 142770 116006 142822 116058
rect 142874 116006 142926 116058
rect 142978 116006 173438 116058
rect 173490 116006 173542 116058
rect 173594 116006 173646 116058
rect 173698 116006 178640 116058
rect 1344 115972 178640 116006
rect 4398 115890 4450 115902
rect 4398 115826 4450 115838
rect 7534 115890 7586 115902
rect 7534 115826 7586 115838
rect 21758 115890 21810 115902
rect 21758 115826 21810 115838
rect 26462 115890 26514 115902
rect 26462 115826 26514 115838
rect 31166 115890 31218 115902
rect 31166 115826 31218 115838
rect 31614 115890 31666 115902
rect 31614 115826 31666 115838
rect 45278 115890 45330 115902
rect 45278 115826 45330 115838
rect 49982 115890 50034 115902
rect 49982 115826 50034 115838
rect 54686 115890 54738 115902
rect 54686 115826 54738 115838
rect 68798 115890 68850 115902
rect 68798 115826 68850 115838
rect 73726 115890 73778 115902
rect 73726 115826 73778 115838
rect 78206 115890 78258 115902
rect 78206 115826 78258 115838
rect 78654 115890 78706 115902
rect 78654 115826 78706 115838
rect 92318 115890 92370 115902
rect 92318 115826 92370 115838
rect 97246 115890 97298 115902
rect 97246 115826 97298 115838
rect 101726 115890 101778 115902
rect 101726 115826 101778 115838
rect 106318 115890 106370 115902
rect 106318 115826 106370 115838
rect 111134 115890 111186 115902
rect 111134 115826 111186 115838
rect 115838 115890 115890 115902
rect 115838 115826 115890 115838
rect 121102 115890 121154 115902
rect 121102 115826 121154 115838
rect 125134 115890 125186 115902
rect 125134 115826 125186 115838
rect 126926 115890 126978 115902
rect 126926 115826 126978 115838
rect 129838 115890 129890 115902
rect 129838 115826 129890 115838
rect 134654 115890 134706 115902
rect 134654 115826 134706 115838
rect 139358 115890 139410 115902
rect 139358 115826 139410 115838
rect 144062 115890 144114 115902
rect 144062 115826 144114 115838
rect 148766 115890 148818 115902
rect 148766 115826 148818 115838
rect 150446 115890 150498 115902
rect 150446 115826 150498 115838
rect 153470 115890 153522 115902
rect 153470 115826 153522 115838
rect 155262 115890 155314 115902
rect 155262 115826 155314 115838
rect 158174 115890 158226 115902
rect 158174 115826 158226 115838
rect 162878 115890 162930 115902
rect 162878 115826 162930 115838
rect 167582 115890 167634 115902
rect 167582 115826 167634 115838
rect 170942 115890 170994 115902
rect 170942 115826 170994 115838
rect 178110 115890 178162 115902
rect 178110 115826 178162 115838
rect 12014 115778 12066 115790
rect 12014 115714 12066 115726
rect 16942 115778 16994 115790
rect 35534 115778 35586 115790
rect 18610 115726 18622 115778
rect 18674 115726 18686 115778
rect 16942 115714 16994 115726
rect 35534 115714 35586 115726
rect 40574 115778 40626 115790
rect 40574 115714 40626 115726
rect 55134 115778 55186 115790
rect 55134 115714 55186 115726
rect 59054 115778 59106 115790
rect 59054 115714 59106 115726
rect 64094 115778 64146 115790
rect 64094 115714 64146 115726
rect 82574 115778 82626 115790
rect 94434 115726 94446 115778
rect 94498 115726 94510 115778
rect 108546 115726 108558 115778
rect 108610 115726 108622 115778
rect 118514 115726 118526 115778
rect 118578 115726 118590 115778
rect 132626 115726 132638 115778
rect 132690 115726 132702 115778
rect 142034 115726 142046 115778
rect 142098 115726 142110 115778
rect 82574 115714 82626 115726
rect 4734 115666 4786 115678
rect 4734 115602 4786 115614
rect 5182 115666 5234 115678
rect 5182 115602 5234 115614
rect 7198 115666 7250 115678
rect 7198 115602 7250 115614
rect 7982 115666 8034 115678
rect 7982 115602 8034 115614
rect 11118 115666 11170 115678
rect 11118 115602 11170 115614
rect 11678 115666 11730 115678
rect 16046 115666 16098 115678
rect 20862 115666 20914 115678
rect 25566 115666 25618 115678
rect 30270 115666 30322 115678
rect 34638 115666 34690 115678
rect 12562 115614 12574 115666
rect 12626 115614 12638 115666
rect 16706 115614 16718 115666
rect 16770 115614 16782 115666
rect 17714 115614 17726 115666
rect 17778 115614 17790 115666
rect 21522 115614 21534 115666
rect 21586 115614 21598 115666
rect 26226 115614 26238 115666
rect 26290 115614 26302 115666
rect 30930 115614 30942 115666
rect 30994 115614 31006 115666
rect 11678 115602 11730 115614
rect 16046 115602 16098 115614
rect 20862 115602 20914 115614
rect 25566 115602 25618 115614
rect 30270 115602 30322 115614
rect 34638 115602 34690 115614
rect 35198 115666 35250 115678
rect 39678 115666 39730 115678
rect 36082 115614 36094 115666
rect 36146 115614 36158 115666
rect 35198 115602 35250 115614
rect 39678 115602 39730 115614
rect 40238 115666 40290 115678
rect 44382 115666 44434 115678
rect 48750 115666 48802 115678
rect 58718 115666 58770 115678
rect 63758 115666 63810 115678
rect 82238 115666 82290 115678
rect 91982 115666 92034 115678
rect 96462 115666 96514 115678
rect 41570 115614 41582 115666
rect 41634 115614 41646 115666
rect 45042 115614 45054 115666
rect 45106 115614 45118 115666
rect 49746 115614 49758 115666
rect 49810 115614 49822 115666
rect 54450 115614 54462 115666
rect 54514 115614 54526 115666
rect 59602 115614 59614 115666
rect 59666 115614 59678 115666
rect 68562 115614 68574 115666
rect 68626 115614 68638 115666
rect 73490 115614 73502 115666
rect 73554 115614 73566 115666
rect 77970 115614 77982 115666
rect 78034 115614 78046 115666
rect 83122 115614 83134 115666
rect 83186 115614 83198 115666
rect 87266 115614 87278 115666
rect 87330 115614 87342 115666
rect 95330 115614 95342 115666
rect 95394 115614 95406 115666
rect 40238 115602 40290 115614
rect 44382 115602 44434 115614
rect 48750 115602 48802 115614
rect 58718 115602 58770 115614
rect 63758 115602 63810 115614
rect 82238 115602 82290 115614
rect 91982 115602 92034 115614
rect 96462 115602 96514 115614
rect 97582 115666 97634 115678
rect 97582 115602 97634 115614
rect 100830 115666 100882 115678
rect 100830 115602 100882 115614
rect 101390 115666 101442 115678
rect 101390 115602 101442 115614
rect 105422 115666 105474 115678
rect 105422 115602 105474 115614
rect 105982 115666 106034 115678
rect 110798 115666 110850 115678
rect 109218 115614 109230 115666
rect 109282 115614 109294 115666
rect 105982 115602 106034 115614
rect 110798 115602 110850 115614
rect 114942 115666 114994 115678
rect 114942 115602 114994 115614
rect 115502 115666 115554 115678
rect 120318 115666 120370 115678
rect 124238 115666 124290 115678
rect 117618 115614 117630 115666
rect 117682 115614 117694 115666
rect 121314 115614 121326 115666
rect 121378 115614 121390 115666
rect 115502 115602 115554 115614
rect 120318 115602 120370 115614
rect 124238 115602 124290 115614
rect 124798 115666 124850 115678
rect 124798 115602 124850 115614
rect 128942 115666 128994 115678
rect 133758 115666 133810 115678
rect 129602 115614 129614 115666
rect 129666 115614 129678 115666
rect 131730 115614 131742 115666
rect 131794 115614 131806 115666
rect 128942 115602 128994 115614
rect 133758 115602 133810 115614
rect 134318 115666 134370 115678
rect 134318 115602 134370 115614
rect 138462 115666 138514 115678
rect 143166 115666 143218 115678
rect 147870 115666 147922 115678
rect 152126 115666 152178 115678
rect 157278 115666 157330 115678
rect 139122 115614 139134 115666
rect 139186 115614 139198 115666
rect 141138 115614 141150 115666
rect 141202 115614 141214 115666
rect 143826 115614 143838 115666
rect 143890 115614 143902 115666
rect 148530 115614 148542 115666
rect 148594 115614 148606 115666
rect 153234 115614 153246 115666
rect 153298 115614 153310 115666
rect 138462 115602 138514 115614
rect 143166 115602 143218 115614
rect 147870 115602 147922 115614
rect 152126 115602 152178 115614
rect 157278 115602 157330 115614
rect 157838 115666 157890 115678
rect 157838 115602 157890 115614
rect 161982 115666 162034 115678
rect 161982 115602 162034 115614
rect 162542 115666 162594 115678
rect 162542 115602 162594 115614
rect 166686 115666 166738 115678
rect 166686 115602 166738 115614
rect 167246 115666 167298 115678
rect 167246 115602 167298 115614
rect 170046 115666 170098 115678
rect 170046 115602 170098 115614
rect 170606 115666 170658 115678
rect 170606 115602 170658 115614
rect 6638 115554 6690 115566
rect 53790 115554 53842 115566
rect 13234 115502 13246 115554
rect 13298 115502 13310 115554
rect 36754 115502 36766 115554
rect 36818 115502 36830 115554
rect 42242 115502 42254 115554
rect 42306 115502 42318 115554
rect 6638 115490 6690 115502
rect 53790 115490 53842 115502
rect 58158 115554 58210 115566
rect 63198 115554 63250 115566
rect 60274 115502 60286 115554
rect 60338 115502 60350 115554
rect 58158 115490 58210 115502
rect 63198 115490 63250 115502
rect 67902 115554 67954 115566
rect 67902 115490 67954 115502
rect 72606 115554 72658 115566
rect 72606 115490 72658 115502
rect 77310 115554 77362 115566
rect 77310 115490 77362 115502
rect 81678 115554 81730 115566
rect 91422 115554 91474 115566
rect 83794 115502 83806 115554
rect 83858 115502 83870 115554
rect 87938 115502 87950 115554
rect 88002 115502 88014 115554
rect 81678 115490 81730 115502
rect 91422 115490 91474 115502
rect 95902 115554 95954 115566
rect 95902 115490 95954 115502
rect 102174 115554 102226 115566
rect 102174 115490 102226 115502
rect 110014 115554 110066 115566
rect 110014 115490 110066 115502
rect 113038 115554 113090 115566
rect 113038 115490 113090 115502
rect 117182 115554 117234 115566
rect 117182 115490 117234 115502
rect 131294 115554 131346 115566
rect 131294 115490 131346 115502
rect 136894 115554 136946 115566
rect 136894 115490 136946 115502
rect 140702 115554 140754 115566
rect 140702 115490 140754 115502
rect 1344 115274 178640 115308
rect 1344 115222 4478 115274
rect 4530 115222 4582 115274
rect 4634 115222 4686 115274
rect 4738 115222 35198 115274
rect 35250 115222 35302 115274
rect 35354 115222 35406 115274
rect 35458 115222 65918 115274
rect 65970 115222 66022 115274
rect 66074 115222 66126 115274
rect 66178 115222 96638 115274
rect 96690 115222 96742 115274
rect 96794 115222 96846 115274
rect 96898 115222 127358 115274
rect 127410 115222 127462 115274
rect 127514 115222 127566 115274
rect 127618 115222 158078 115274
rect 158130 115222 158182 115274
rect 158234 115222 158286 115274
rect 158338 115222 178640 115274
rect 1344 115188 178640 115222
rect 110462 114994 110514 115006
rect 64978 114942 64990 114994
rect 65042 114942 65054 114994
rect 110462 114930 110514 114942
rect 86718 114882 86770 114894
rect 64306 114830 64318 114882
rect 64370 114830 64382 114882
rect 86718 114818 86770 114830
rect 87614 114882 87666 114894
rect 87614 114818 87666 114830
rect 87278 114770 87330 114782
rect 87278 114706 87330 114718
rect 1344 114490 178640 114524
rect 1344 114438 19838 114490
rect 19890 114438 19942 114490
rect 19994 114438 20046 114490
rect 20098 114438 50558 114490
rect 50610 114438 50662 114490
rect 50714 114438 50766 114490
rect 50818 114438 81278 114490
rect 81330 114438 81382 114490
rect 81434 114438 81486 114490
rect 81538 114438 111998 114490
rect 112050 114438 112102 114490
rect 112154 114438 112206 114490
rect 112258 114438 142718 114490
rect 142770 114438 142822 114490
rect 142874 114438 142926 114490
rect 142978 114438 173438 114490
rect 173490 114438 173542 114490
rect 173594 114438 173646 114490
rect 173698 114438 178640 114490
rect 1344 114404 178640 114438
rect 1344 113706 178640 113740
rect 1344 113654 4478 113706
rect 4530 113654 4582 113706
rect 4634 113654 4686 113706
rect 4738 113654 35198 113706
rect 35250 113654 35302 113706
rect 35354 113654 35406 113706
rect 35458 113654 65918 113706
rect 65970 113654 66022 113706
rect 66074 113654 66126 113706
rect 66178 113654 96638 113706
rect 96690 113654 96742 113706
rect 96794 113654 96846 113706
rect 96898 113654 127358 113706
rect 127410 113654 127462 113706
rect 127514 113654 127566 113706
rect 127618 113654 158078 113706
rect 158130 113654 158182 113706
rect 158234 113654 158286 113706
rect 158338 113654 178640 113706
rect 1344 113620 178640 113654
rect 1344 112922 178640 112956
rect 1344 112870 19838 112922
rect 19890 112870 19942 112922
rect 19994 112870 20046 112922
rect 20098 112870 50558 112922
rect 50610 112870 50662 112922
rect 50714 112870 50766 112922
rect 50818 112870 81278 112922
rect 81330 112870 81382 112922
rect 81434 112870 81486 112922
rect 81538 112870 111998 112922
rect 112050 112870 112102 112922
rect 112154 112870 112206 112922
rect 112258 112870 142718 112922
rect 142770 112870 142822 112922
rect 142874 112870 142926 112922
rect 142978 112870 173438 112922
rect 173490 112870 173542 112922
rect 173594 112870 173646 112922
rect 173698 112870 178640 112922
rect 1344 112836 178640 112870
rect 1344 112138 178640 112172
rect 1344 112086 4478 112138
rect 4530 112086 4582 112138
rect 4634 112086 4686 112138
rect 4738 112086 35198 112138
rect 35250 112086 35302 112138
rect 35354 112086 35406 112138
rect 35458 112086 65918 112138
rect 65970 112086 66022 112138
rect 66074 112086 66126 112138
rect 66178 112086 96638 112138
rect 96690 112086 96742 112138
rect 96794 112086 96846 112138
rect 96898 112086 127358 112138
rect 127410 112086 127462 112138
rect 127514 112086 127566 112138
rect 127618 112086 158078 112138
rect 158130 112086 158182 112138
rect 158234 112086 158286 112138
rect 158338 112086 178640 112138
rect 1344 112052 178640 112086
rect 1344 111354 178640 111388
rect 1344 111302 19838 111354
rect 19890 111302 19942 111354
rect 19994 111302 20046 111354
rect 20098 111302 50558 111354
rect 50610 111302 50662 111354
rect 50714 111302 50766 111354
rect 50818 111302 81278 111354
rect 81330 111302 81382 111354
rect 81434 111302 81486 111354
rect 81538 111302 111998 111354
rect 112050 111302 112102 111354
rect 112154 111302 112206 111354
rect 112258 111302 142718 111354
rect 142770 111302 142822 111354
rect 142874 111302 142926 111354
rect 142978 111302 173438 111354
rect 173490 111302 173542 111354
rect 173594 111302 173646 111354
rect 173698 111302 178640 111354
rect 1344 111268 178640 111302
rect 1344 110570 178640 110604
rect 1344 110518 4478 110570
rect 4530 110518 4582 110570
rect 4634 110518 4686 110570
rect 4738 110518 35198 110570
rect 35250 110518 35302 110570
rect 35354 110518 35406 110570
rect 35458 110518 65918 110570
rect 65970 110518 66022 110570
rect 66074 110518 66126 110570
rect 66178 110518 96638 110570
rect 96690 110518 96742 110570
rect 96794 110518 96846 110570
rect 96898 110518 127358 110570
rect 127410 110518 127462 110570
rect 127514 110518 127566 110570
rect 127618 110518 158078 110570
rect 158130 110518 158182 110570
rect 158234 110518 158286 110570
rect 158338 110518 178640 110570
rect 1344 110484 178640 110518
rect 1344 109786 178640 109820
rect 1344 109734 19838 109786
rect 19890 109734 19942 109786
rect 19994 109734 20046 109786
rect 20098 109734 50558 109786
rect 50610 109734 50662 109786
rect 50714 109734 50766 109786
rect 50818 109734 81278 109786
rect 81330 109734 81382 109786
rect 81434 109734 81486 109786
rect 81538 109734 111998 109786
rect 112050 109734 112102 109786
rect 112154 109734 112206 109786
rect 112258 109734 142718 109786
rect 142770 109734 142822 109786
rect 142874 109734 142926 109786
rect 142978 109734 173438 109786
rect 173490 109734 173542 109786
rect 173594 109734 173646 109786
rect 173698 109734 178640 109786
rect 1344 109700 178640 109734
rect 1344 109002 178640 109036
rect 1344 108950 4478 109002
rect 4530 108950 4582 109002
rect 4634 108950 4686 109002
rect 4738 108950 35198 109002
rect 35250 108950 35302 109002
rect 35354 108950 35406 109002
rect 35458 108950 65918 109002
rect 65970 108950 66022 109002
rect 66074 108950 66126 109002
rect 66178 108950 96638 109002
rect 96690 108950 96742 109002
rect 96794 108950 96846 109002
rect 96898 108950 127358 109002
rect 127410 108950 127462 109002
rect 127514 108950 127566 109002
rect 127618 108950 158078 109002
rect 158130 108950 158182 109002
rect 158234 108950 158286 109002
rect 158338 108950 178640 109002
rect 1344 108916 178640 108950
rect 1344 108218 178640 108252
rect 1344 108166 19838 108218
rect 19890 108166 19942 108218
rect 19994 108166 20046 108218
rect 20098 108166 50558 108218
rect 50610 108166 50662 108218
rect 50714 108166 50766 108218
rect 50818 108166 81278 108218
rect 81330 108166 81382 108218
rect 81434 108166 81486 108218
rect 81538 108166 111998 108218
rect 112050 108166 112102 108218
rect 112154 108166 112206 108218
rect 112258 108166 142718 108218
rect 142770 108166 142822 108218
rect 142874 108166 142926 108218
rect 142978 108166 173438 108218
rect 173490 108166 173542 108218
rect 173594 108166 173646 108218
rect 173698 108166 178640 108218
rect 1344 108132 178640 108166
rect 1344 107434 178640 107468
rect 1344 107382 4478 107434
rect 4530 107382 4582 107434
rect 4634 107382 4686 107434
rect 4738 107382 35198 107434
rect 35250 107382 35302 107434
rect 35354 107382 35406 107434
rect 35458 107382 65918 107434
rect 65970 107382 66022 107434
rect 66074 107382 66126 107434
rect 66178 107382 96638 107434
rect 96690 107382 96742 107434
rect 96794 107382 96846 107434
rect 96898 107382 127358 107434
rect 127410 107382 127462 107434
rect 127514 107382 127566 107434
rect 127618 107382 158078 107434
rect 158130 107382 158182 107434
rect 158234 107382 158286 107434
rect 158338 107382 178640 107434
rect 1344 107348 178640 107382
rect 1344 106650 178640 106684
rect 1344 106598 19838 106650
rect 19890 106598 19942 106650
rect 19994 106598 20046 106650
rect 20098 106598 50558 106650
rect 50610 106598 50662 106650
rect 50714 106598 50766 106650
rect 50818 106598 81278 106650
rect 81330 106598 81382 106650
rect 81434 106598 81486 106650
rect 81538 106598 111998 106650
rect 112050 106598 112102 106650
rect 112154 106598 112206 106650
rect 112258 106598 142718 106650
rect 142770 106598 142822 106650
rect 142874 106598 142926 106650
rect 142978 106598 173438 106650
rect 173490 106598 173542 106650
rect 173594 106598 173646 106650
rect 173698 106598 178640 106650
rect 1344 106564 178640 106598
rect 1344 105866 178640 105900
rect 1344 105814 4478 105866
rect 4530 105814 4582 105866
rect 4634 105814 4686 105866
rect 4738 105814 35198 105866
rect 35250 105814 35302 105866
rect 35354 105814 35406 105866
rect 35458 105814 65918 105866
rect 65970 105814 66022 105866
rect 66074 105814 66126 105866
rect 66178 105814 96638 105866
rect 96690 105814 96742 105866
rect 96794 105814 96846 105866
rect 96898 105814 127358 105866
rect 127410 105814 127462 105866
rect 127514 105814 127566 105866
rect 127618 105814 158078 105866
rect 158130 105814 158182 105866
rect 158234 105814 158286 105866
rect 158338 105814 178640 105866
rect 1344 105780 178640 105814
rect 1344 105082 178640 105116
rect 1344 105030 19838 105082
rect 19890 105030 19942 105082
rect 19994 105030 20046 105082
rect 20098 105030 50558 105082
rect 50610 105030 50662 105082
rect 50714 105030 50766 105082
rect 50818 105030 81278 105082
rect 81330 105030 81382 105082
rect 81434 105030 81486 105082
rect 81538 105030 111998 105082
rect 112050 105030 112102 105082
rect 112154 105030 112206 105082
rect 112258 105030 142718 105082
rect 142770 105030 142822 105082
rect 142874 105030 142926 105082
rect 142978 105030 173438 105082
rect 173490 105030 173542 105082
rect 173594 105030 173646 105082
rect 173698 105030 178640 105082
rect 1344 104996 178640 105030
rect 1344 104298 178640 104332
rect 1344 104246 4478 104298
rect 4530 104246 4582 104298
rect 4634 104246 4686 104298
rect 4738 104246 35198 104298
rect 35250 104246 35302 104298
rect 35354 104246 35406 104298
rect 35458 104246 65918 104298
rect 65970 104246 66022 104298
rect 66074 104246 66126 104298
rect 66178 104246 96638 104298
rect 96690 104246 96742 104298
rect 96794 104246 96846 104298
rect 96898 104246 127358 104298
rect 127410 104246 127462 104298
rect 127514 104246 127566 104298
rect 127618 104246 158078 104298
rect 158130 104246 158182 104298
rect 158234 104246 158286 104298
rect 158338 104246 178640 104298
rect 1344 104212 178640 104246
rect 1344 103514 178640 103548
rect 1344 103462 19838 103514
rect 19890 103462 19942 103514
rect 19994 103462 20046 103514
rect 20098 103462 50558 103514
rect 50610 103462 50662 103514
rect 50714 103462 50766 103514
rect 50818 103462 81278 103514
rect 81330 103462 81382 103514
rect 81434 103462 81486 103514
rect 81538 103462 111998 103514
rect 112050 103462 112102 103514
rect 112154 103462 112206 103514
rect 112258 103462 142718 103514
rect 142770 103462 142822 103514
rect 142874 103462 142926 103514
rect 142978 103462 173438 103514
rect 173490 103462 173542 103514
rect 173594 103462 173646 103514
rect 173698 103462 178640 103514
rect 1344 103428 178640 103462
rect 1344 102730 178640 102764
rect 1344 102678 4478 102730
rect 4530 102678 4582 102730
rect 4634 102678 4686 102730
rect 4738 102678 35198 102730
rect 35250 102678 35302 102730
rect 35354 102678 35406 102730
rect 35458 102678 65918 102730
rect 65970 102678 66022 102730
rect 66074 102678 66126 102730
rect 66178 102678 96638 102730
rect 96690 102678 96742 102730
rect 96794 102678 96846 102730
rect 96898 102678 127358 102730
rect 127410 102678 127462 102730
rect 127514 102678 127566 102730
rect 127618 102678 158078 102730
rect 158130 102678 158182 102730
rect 158234 102678 158286 102730
rect 158338 102678 178640 102730
rect 1344 102644 178640 102678
rect 1344 101946 178640 101980
rect 1344 101894 19838 101946
rect 19890 101894 19942 101946
rect 19994 101894 20046 101946
rect 20098 101894 50558 101946
rect 50610 101894 50662 101946
rect 50714 101894 50766 101946
rect 50818 101894 81278 101946
rect 81330 101894 81382 101946
rect 81434 101894 81486 101946
rect 81538 101894 111998 101946
rect 112050 101894 112102 101946
rect 112154 101894 112206 101946
rect 112258 101894 142718 101946
rect 142770 101894 142822 101946
rect 142874 101894 142926 101946
rect 142978 101894 173438 101946
rect 173490 101894 173542 101946
rect 173594 101894 173646 101946
rect 173698 101894 178640 101946
rect 1344 101860 178640 101894
rect 1344 101162 178640 101196
rect 1344 101110 4478 101162
rect 4530 101110 4582 101162
rect 4634 101110 4686 101162
rect 4738 101110 35198 101162
rect 35250 101110 35302 101162
rect 35354 101110 35406 101162
rect 35458 101110 65918 101162
rect 65970 101110 66022 101162
rect 66074 101110 66126 101162
rect 66178 101110 96638 101162
rect 96690 101110 96742 101162
rect 96794 101110 96846 101162
rect 96898 101110 127358 101162
rect 127410 101110 127462 101162
rect 127514 101110 127566 101162
rect 127618 101110 158078 101162
rect 158130 101110 158182 101162
rect 158234 101110 158286 101162
rect 158338 101110 178640 101162
rect 1344 101076 178640 101110
rect 1344 100378 178640 100412
rect 1344 100326 19838 100378
rect 19890 100326 19942 100378
rect 19994 100326 20046 100378
rect 20098 100326 50558 100378
rect 50610 100326 50662 100378
rect 50714 100326 50766 100378
rect 50818 100326 81278 100378
rect 81330 100326 81382 100378
rect 81434 100326 81486 100378
rect 81538 100326 111998 100378
rect 112050 100326 112102 100378
rect 112154 100326 112206 100378
rect 112258 100326 142718 100378
rect 142770 100326 142822 100378
rect 142874 100326 142926 100378
rect 142978 100326 173438 100378
rect 173490 100326 173542 100378
rect 173594 100326 173646 100378
rect 173698 100326 178640 100378
rect 1344 100292 178640 100326
rect 1344 99594 178640 99628
rect 1344 99542 4478 99594
rect 4530 99542 4582 99594
rect 4634 99542 4686 99594
rect 4738 99542 35198 99594
rect 35250 99542 35302 99594
rect 35354 99542 35406 99594
rect 35458 99542 65918 99594
rect 65970 99542 66022 99594
rect 66074 99542 66126 99594
rect 66178 99542 96638 99594
rect 96690 99542 96742 99594
rect 96794 99542 96846 99594
rect 96898 99542 127358 99594
rect 127410 99542 127462 99594
rect 127514 99542 127566 99594
rect 127618 99542 158078 99594
rect 158130 99542 158182 99594
rect 158234 99542 158286 99594
rect 158338 99542 178640 99594
rect 1344 99508 178640 99542
rect 1344 98810 178640 98844
rect 1344 98758 19838 98810
rect 19890 98758 19942 98810
rect 19994 98758 20046 98810
rect 20098 98758 50558 98810
rect 50610 98758 50662 98810
rect 50714 98758 50766 98810
rect 50818 98758 81278 98810
rect 81330 98758 81382 98810
rect 81434 98758 81486 98810
rect 81538 98758 111998 98810
rect 112050 98758 112102 98810
rect 112154 98758 112206 98810
rect 112258 98758 142718 98810
rect 142770 98758 142822 98810
rect 142874 98758 142926 98810
rect 142978 98758 173438 98810
rect 173490 98758 173542 98810
rect 173594 98758 173646 98810
rect 173698 98758 178640 98810
rect 1344 98724 178640 98758
rect 1344 98026 178640 98060
rect 1344 97974 4478 98026
rect 4530 97974 4582 98026
rect 4634 97974 4686 98026
rect 4738 97974 35198 98026
rect 35250 97974 35302 98026
rect 35354 97974 35406 98026
rect 35458 97974 65918 98026
rect 65970 97974 66022 98026
rect 66074 97974 66126 98026
rect 66178 97974 96638 98026
rect 96690 97974 96742 98026
rect 96794 97974 96846 98026
rect 96898 97974 127358 98026
rect 127410 97974 127462 98026
rect 127514 97974 127566 98026
rect 127618 97974 158078 98026
rect 158130 97974 158182 98026
rect 158234 97974 158286 98026
rect 158338 97974 178640 98026
rect 1344 97940 178640 97974
rect 1344 97242 178640 97276
rect 1344 97190 19838 97242
rect 19890 97190 19942 97242
rect 19994 97190 20046 97242
rect 20098 97190 50558 97242
rect 50610 97190 50662 97242
rect 50714 97190 50766 97242
rect 50818 97190 81278 97242
rect 81330 97190 81382 97242
rect 81434 97190 81486 97242
rect 81538 97190 111998 97242
rect 112050 97190 112102 97242
rect 112154 97190 112206 97242
rect 112258 97190 142718 97242
rect 142770 97190 142822 97242
rect 142874 97190 142926 97242
rect 142978 97190 173438 97242
rect 173490 97190 173542 97242
rect 173594 97190 173646 97242
rect 173698 97190 178640 97242
rect 1344 97156 178640 97190
rect 1344 96458 178640 96492
rect 1344 96406 4478 96458
rect 4530 96406 4582 96458
rect 4634 96406 4686 96458
rect 4738 96406 35198 96458
rect 35250 96406 35302 96458
rect 35354 96406 35406 96458
rect 35458 96406 65918 96458
rect 65970 96406 66022 96458
rect 66074 96406 66126 96458
rect 66178 96406 96638 96458
rect 96690 96406 96742 96458
rect 96794 96406 96846 96458
rect 96898 96406 127358 96458
rect 127410 96406 127462 96458
rect 127514 96406 127566 96458
rect 127618 96406 158078 96458
rect 158130 96406 158182 96458
rect 158234 96406 158286 96458
rect 158338 96406 178640 96458
rect 1344 96372 178640 96406
rect 1344 95674 178640 95708
rect 1344 95622 19838 95674
rect 19890 95622 19942 95674
rect 19994 95622 20046 95674
rect 20098 95622 50558 95674
rect 50610 95622 50662 95674
rect 50714 95622 50766 95674
rect 50818 95622 81278 95674
rect 81330 95622 81382 95674
rect 81434 95622 81486 95674
rect 81538 95622 111998 95674
rect 112050 95622 112102 95674
rect 112154 95622 112206 95674
rect 112258 95622 142718 95674
rect 142770 95622 142822 95674
rect 142874 95622 142926 95674
rect 142978 95622 173438 95674
rect 173490 95622 173542 95674
rect 173594 95622 173646 95674
rect 173698 95622 178640 95674
rect 1344 95588 178640 95622
rect 1344 94890 178640 94924
rect 1344 94838 4478 94890
rect 4530 94838 4582 94890
rect 4634 94838 4686 94890
rect 4738 94838 35198 94890
rect 35250 94838 35302 94890
rect 35354 94838 35406 94890
rect 35458 94838 65918 94890
rect 65970 94838 66022 94890
rect 66074 94838 66126 94890
rect 66178 94838 96638 94890
rect 96690 94838 96742 94890
rect 96794 94838 96846 94890
rect 96898 94838 127358 94890
rect 127410 94838 127462 94890
rect 127514 94838 127566 94890
rect 127618 94838 158078 94890
rect 158130 94838 158182 94890
rect 158234 94838 158286 94890
rect 158338 94838 178640 94890
rect 1344 94804 178640 94838
rect 1344 94106 178640 94140
rect 1344 94054 19838 94106
rect 19890 94054 19942 94106
rect 19994 94054 20046 94106
rect 20098 94054 50558 94106
rect 50610 94054 50662 94106
rect 50714 94054 50766 94106
rect 50818 94054 81278 94106
rect 81330 94054 81382 94106
rect 81434 94054 81486 94106
rect 81538 94054 111998 94106
rect 112050 94054 112102 94106
rect 112154 94054 112206 94106
rect 112258 94054 142718 94106
rect 142770 94054 142822 94106
rect 142874 94054 142926 94106
rect 142978 94054 173438 94106
rect 173490 94054 173542 94106
rect 173594 94054 173646 94106
rect 173698 94054 178640 94106
rect 1344 94020 178640 94054
rect 1344 93322 178640 93356
rect 1344 93270 4478 93322
rect 4530 93270 4582 93322
rect 4634 93270 4686 93322
rect 4738 93270 35198 93322
rect 35250 93270 35302 93322
rect 35354 93270 35406 93322
rect 35458 93270 65918 93322
rect 65970 93270 66022 93322
rect 66074 93270 66126 93322
rect 66178 93270 96638 93322
rect 96690 93270 96742 93322
rect 96794 93270 96846 93322
rect 96898 93270 127358 93322
rect 127410 93270 127462 93322
rect 127514 93270 127566 93322
rect 127618 93270 158078 93322
rect 158130 93270 158182 93322
rect 158234 93270 158286 93322
rect 158338 93270 178640 93322
rect 1344 93236 178640 93270
rect 1344 92538 178640 92572
rect 1344 92486 19838 92538
rect 19890 92486 19942 92538
rect 19994 92486 20046 92538
rect 20098 92486 50558 92538
rect 50610 92486 50662 92538
rect 50714 92486 50766 92538
rect 50818 92486 81278 92538
rect 81330 92486 81382 92538
rect 81434 92486 81486 92538
rect 81538 92486 111998 92538
rect 112050 92486 112102 92538
rect 112154 92486 112206 92538
rect 112258 92486 142718 92538
rect 142770 92486 142822 92538
rect 142874 92486 142926 92538
rect 142978 92486 173438 92538
rect 173490 92486 173542 92538
rect 173594 92486 173646 92538
rect 173698 92486 178640 92538
rect 1344 92452 178640 92486
rect 1344 91754 178640 91788
rect 1344 91702 4478 91754
rect 4530 91702 4582 91754
rect 4634 91702 4686 91754
rect 4738 91702 35198 91754
rect 35250 91702 35302 91754
rect 35354 91702 35406 91754
rect 35458 91702 65918 91754
rect 65970 91702 66022 91754
rect 66074 91702 66126 91754
rect 66178 91702 96638 91754
rect 96690 91702 96742 91754
rect 96794 91702 96846 91754
rect 96898 91702 127358 91754
rect 127410 91702 127462 91754
rect 127514 91702 127566 91754
rect 127618 91702 158078 91754
rect 158130 91702 158182 91754
rect 158234 91702 158286 91754
rect 158338 91702 178640 91754
rect 1344 91668 178640 91702
rect 1344 90970 178640 91004
rect 1344 90918 19838 90970
rect 19890 90918 19942 90970
rect 19994 90918 20046 90970
rect 20098 90918 50558 90970
rect 50610 90918 50662 90970
rect 50714 90918 50766 90970
rect 50818 90918 81278 90970
rect 81330 90918 81382 90970
rect 81434 90918 81486 90970
rect 81538 90918 111998 90970
rect 112050 90918 112102 90970
rect 112154 90918 112206 90970
rect 112258 90918 142718 90970
rect 142770 90918 142822 90970
rect 142874 90918 142926 90970
rect 142978 90918 173438 90970
rect 173490 90918 173542 90970
rect 173594 90918 173646 90970
rect 173698 90918 178640 90970
rect 1344 90884 178640 90918
rect 1344 90186 178640 90220
rect 1344 90134 4478 90186
rect 4530 90134 4582 90186
rect 4634 90134 4686 90186
rect 4738 90134 35198 90186
rect 35250 90134 35302 90186
rect 35354 90134 35406 90186
rect 35458 90134 65918 90186
rect 65970 90134 66022 90186
rect 66074 90134 66126 90186
rect 66178 90134 96638 90186
rect 96690 90134 96742 90186
rect 96794 90134 96846 90186
rect 96898 90134 127358 90186
rect 127410 90134 127462 90186
rect 127514 90134 127566 90186
rect 127618 90134 158078 90186
rect 158130 90134 158182 90186
rect 158234 90134 158286 90186
rect 158338 90134 178640 90186
rect 1344 90100 178640 90134
rect 1344 89402 178640 89436
rect 1344 89350 19838 89402
rect 19890 89350 19942 89402
rect 19994 89350 20046 89402
rect 20098 89350 50558 89402
rect 50610 89350 50662 89402
rect 50714 89350 50766 89402
rect 50818 89350 81278 89402
rect 81330 89350 81382 89402
rect 81434 89350 81486 89402
rect 81538 89350 111998 89402
rect 112050 89350 112102 89402
rect 112154 89350 112206 89402
rect 112258 89350 142718 89402
rect 142770 89350 142822 89402
rect 142874 89350 142926 89402
rect 142978 89350 173438 89402
rect 173490 89350 173542 89402
rect 173594 89350 173646 89402
rect 173698 89350 178640 89402
rect 1344 89316 178640 89350
rect 1344 88618 178640 88652
rect 1344 88566 4478 88618
rect 4530 88566 4582 88618
rect 4634 88566 4686 88618
rect 4738 88566 35198 88618
rect 35250 88566 35302 88618
rect 35354 88566 35406 88618
rect 35458 88566 65918 88618
rect 65970 88566 66022 88618
rect 66074 88566 66126 88618
rect 66178 88566 96638 88618
rect 96690 88566 96742 88618
rect 96794 88566 96846 88618
rect 96898 88566 127358 88618
rect 127410 88566 127462 88618
rect 127514 88566 127566 88618
rect 127618 88566 158078 88618
rect 158130 88566 158182 88618
rect 158234 88566 158286 88618
rect 158338 88566 178640 88618
rect 1344 88532 178640 88566
rect 1344 87834 178640 87868
rect 1344 87782 19838 87834
rect 19890 87782 19942 87834
rect 19994 87782 20046 87834
rect 20098 87782 50558 87834
rect 50610 87782 50662 87834
rect 50714 87782 50766 87834
rect 50818 87782 81278 87834
rect 81330 87782 81382 87834
rect 81434 87782 81486 87834
rect 81538 87782 111998 87834
rect 112050 87782 112102 87834
rect 112154 87782 112206 87834
rect 112258 87782 142718 87834
rect 142770 87782 142822 87834
rect 142874 87782 142926 87834
rect 142978 87782 173438 87834
rect 173490 87782 173542 87834
rect 173594 87782 173646 87834
rect 173698 87782 178640 87834
rect 1344 87748 178640 87782
rect 1344 87050 178640 87084
rect 1344 86998 4478 87050
rect 4530 86998 4582 87050
rect 4634 86998 4686 87050
rect 4738 86998 35198 87050
rect 35250 86998 35302 87050
rect 35354 86998 35406 87050
rect 35458 86998 65918 87050
rect 65970 86998 66022 87050
rect 66074 86998 66126 87050
rect 66178 86998 96638 87050
rect 96690 86998 96742 87050
rect 96794 86998 96846 87050
rect 96898 86998 127358 87050
rect 127410 86998 127462 87050
rect 127514 86998 127566 87050
rect 127618 86998 158078 87050
rect 158130 86998 158182 87050
rect 158234 86998 158286 87050
rect 158338 86998 178640 87050
rect 1344 86964 178640 86998
rect 1344 86266 178640 86300
rect 1344 86214 19838 86266
rect 19890 86214 19942 86266
rect 19994 86214 20046 86266
rect 20098 86214 50558 86266
rect 50610 86214 50662 86266
rect 50714 86214 50766 86266
rect 50818 86214 81278 86266
rect 81330 86214 81382 86266
rect 81434 86214 81486 86266
rect 81538 86214 111998 86266
rect 112050 86214 112102 86266
rect 112154 86214 112206 86266
rect 112258 86214 142718 86266
rect 142770 86214 142822 86266
rect 142874 86214 142926 86266
rect 142978 86214 173438 86266
rect 173490 86214 173542 86266
rect 173594 86214 173646 86266
rect 173698 86214 178640 86266
rect 1344 86180 178640 86214
rect 1344 85482 178640 85516
rect 1344 85430 4478 85482
rect 4530 85430 4582 85482
rect 4634 85430 4686 85482
rect 4738 85430 35198 85482
rect 35250 85430 35302 85482
rect 35354 85430 35406 85482
rect 35458 85430 65918 85482
rect 65970 85430 66022 85482
rect 66074 85430 66126 85482
rect 66178 85430 96638 85482
rect 96690 85430 96742 85482
rect 96794 85430 96846 85482
rect 96898 85430 127358 85482
rect 127410 85430 127462 85482
rect 127514 85430 127566 85482
rect 127618 85430 158078 85482
rect 158130 85430 158182 85482
rect 158234 85430 158286 85482
rect 158338 85430 178640 85482
rect 1344 85396 178640 85430
rect 1344 84698 178640 84732
rect 1344 84646 19838 84698
rect 19890 84646 19942 84698
rect 19994 84646 20046 84698
rect 20098 84646 50558 84698
rect 50610 84646 50662 84698
rect 50714 84646 50766 84698
rect 50818 84646 81278 84698
rect 81330 84646 81382 84698
rect 81434 84646 81486 84698
rect 81538 84646 111998 84698
rect 112050 84646 112102 84698
rect 112154 84646 112206 84698
rect 112258 84646 142718 84698
rect 142770 84646 142822 84698
rect 142874 84646 142926 84698
rect 142978 84646 173438 84698
rect 173490 84646 173542 84698
rect 173594 84646 173646 84698
rect 173698 84646 178640 84698
rect 1344 84612 178640 84646
rect 1344 83914 178640 83948
rect 1344 83862 4478 83914
rect 4530 83862 4582 83914
rect 4634 83862 4686 83914
rect 4738 83862 35198 83914
rect 35250 83862 35302 83914
rect 35354 83862 35406 83914
rect 35458 83862 65918 83914
rect 65970 83862 66022 83914
rect 66074 83862 66126 83914
rect 66178 83862 96638 83914
rect 96690 83862 96742 83914
rect 96794 83862 96846 83914
rect 96898 83862 127358 83914
rect 127410 83862 127462 83914
rect 127514 83862 127566 83914
rect 127618 83862 158078 83914
rect 158130 83862 158182 83914
rect 158234 83862 158286 83914
rect 158338 83862 178640 83914
rect 1344 83828 178640 83862
rect 1344 83130 178640 83164
rect 1344 83078 19838 83130
rect 19890 83078 19942 83130
rect 19994 83078 20046 83130
rect 20098 83078 50558 83130
rect 50610 83078 50662 83130
rect 50714 83078 50766 83130
rect 50818 83078 81278 83130
rect 81330 83078 81382 83130
rect 81434 83078 81486 83130
rect 81538 83078 111998 83130
rect 112050 83078 112102 83130
rect 112154 83078 112206 83130
rect 112258 83078 142718 83130
rect 142770 83078 142822 83130
rect 142874 83078 142926 83130
rect 142978 83078 173438 83130
rect 173490 83078 173542 83130
rect 173594 83078 173646 83130
rect 173698 83078 178640 83130
rect 1344 83044 178640 83078
rect 1344 82346 178640 82380
rect 1344 82294 4478 82346
rect 4530 82294 4582 82346
rect 4634 82294 4686 82346
rect 4738 82294 35198 82346
rect 35250 82294 35302 82346
rect 35354 82294 35406 82346
rect 35458 82294 65918 82346
rect 65970 82294 66022 82346
rect 66074 82294 66126 82346
rect 66178 82294 96638 82346
rect 96690 82294 96742 82346
rect 96794 82294 96846 82346
rect 96898 82294 127358 82346
rect 127410 82294 127462 82346
rect 127514 82294 127566 82346
rect 127618 82294 158078 82346
rect 158130 82294 158182 82346
rect 158234 82294 158286 82346
rect 158338 82294 178640 82346
rect 1344 82260 178640 82294
rect 1344 81562 178640 81596
rect 1344 81510 19838 81562
rect 19890 81510 19942 81562
rect 19994 81510 20046 81562
rect 20098 81510 50558 81562
rect 50610 81510 50662 81562
rect 50714 81510 50766 81562
rect 50818 81510 81278 81562
rect 81330 81510 81382 81562
rect 81434 81510 81486 81562
rect 81538 81510 111998 81562
rect 112050 81510 112102 81562
rect 112154 81510 112206 81562
rect 112258 81510 142718 81562
rect 142770 81510 142822 81562
rect 142874 81510 142926 81562
rect 142978 81510 173438 81562
rect 173490 81510 173542 81562
rect 173594 81510 173646 81562
rect 173698 81510 178640 81562
rect 1344 81476 178640 81510
rect 1344 80778 178640 80812
rect 1344 80726 4478 80778
rect 4530 80726 4582 80778
rect 4634 80726 4686 80778
rect 4738 80726 35198 80778
rect 35250 80726 35302 80778
rect 35354 80726 35406 80778
rect 35458 80726 65918 80778
rect 65970 80726 66022 80778
rect 66074 80726 66126 80778
rect 66178 80726 96638 80778
rect 96690 80726 96742 80778
rect 96794 80726 96846 80778
rect 96898 80726 127358 80778
rect 127410 80726 127462 80778
rect 127514 80726 127566 80778
rect 127618 80726 158078 80778
rect 158130 80726 158182 80778
rect 158234 80726 158286 80778
rect 158338 80726 178640 80778
rect 1344 80692 178640 80726
rect 1344 79994 178640 80028
rect 1344 79942 19838 79994
rect 19890 79942 19942 79994
rect 19994 79942 20046 79994
rect 20098 79942 50558 79994
rect 50610 79942 50662 79994
rect 50714 79942 50766 79994
rect 50818 79942 81278 79994
rect 81330 79942 81382 79994
rect 81434 79942 81486 79994
rect 81538 79942 111998 79994
rect 112050 79942 112102 79994
rect 112154 79942 112206 79994
rect 112258 79942 142718 79994
rect 142770 79942 142822 79994
rect 142874 79942 142926 79994
rect 142978 79942 173438 79994
rect 173490 79942 173542 79994
rect 173594 79942 173646 79994
rect 173698 79942 178640 79994
rect 1344 79908 178640 79942
rect 1344 79210 178640 79244
rect 1344 79158 4478 79210
rect 4530 79158 4582 79210
rect 4634 79158 4686 79210
rect 4738 79158 35198 79210
rect 35250 79158 35302 79210
rect 35354 79158 35406 79210
rect 35458 79158 65918 79210
rect 65970 79158 66022 79210
rect 66074 79158 66126 79210
rect 66178 79158 96638 79210
rect 96690 79158 96742 79210
rect 96794 79158 96846 79210
rect 96898 79158 127358 79210
rect 127410 79158 127462 79210
rect 127514 79158 127566 79210
rect 127618 79158 158078 79210
rect 158130 79158 158182 79210
rect 158234 79158 158286 79210
rect 158338 79158 178640 79210
rect 1344 79124 178640 79158
rect 1344 78426 178640 78460
rect 1344 78374 19838 78426
rect 19890 78374 19942 78426
rect 19994 78374 20046 78426
rect 20098 78374 50558 78426
rect 50610 78374 50662 78426
rect 50714 78374 50766 78426
rect 50818 78374 81278 78426
rect 81330 78374 81382 78426
rect 81434 78374 81486 78426
rect 81538 78374 111998 78426
rect 112050 78374 112102 78426
rect 112154 78374 112206 78426
rect 112258 78374 142718 78426
rect 142770 78374 142822 78426
rect 142874 78374 142926 78426
rect 142978 78374 173438 78426
rect 173490 78374 173542 78426
rect 173594 78374 173646 78426
rect 173698 78374 178640 78426
rect 1344 78340 178640 78374
rect 1344 77642 178640 77676
rect 1344 77590 4478 77642
rect 4530 77590 4582 77642
rect 4634 77590 4686 77642
rect 4738 77590 35198 77642
rect 35250 77590 35302 77642
rect 35354 77590 35406 77642
rect 35458 77590 65918 77642
rect 65970 77590 66022 77642
rect 66074 77590 66126 77642
rect 66178 77590 96638 77642
rect 96690 77590 96742 77642
rect 96794 77590 96846 77642
rect 96898 77590 127358 77642
rect 127410 77590 127462 77642
rect 127514 77590 127566 77642
rect 127618 77590 158078 77642
rect 158130 77590 158182 77642
rect 158234 77590 158286 77642
rect 158338 77590 178640 77642
rect 1344 77556 178640 77590
rect 1344 76858 178640 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 81278 76858
rect 81330 76806 81382 76858
rect 81434 76806 81486 76858
rect 81538 76806 111998 76858
rect 112050 76806 112102 76858
rect 112154 76806 112206 76858
rect 112258 76806 142718 76858
rect 142770 76806 142822 76858
rect 142874 76806 142926 76858
rect 142978 76806 173438 76858
rect 173490 76806 173542 76858
rect 173594 76806 173646 76858
rect 173698 76806 178640 76858
rect 1344 76772 178640 76806
rect 1344 76074 178640 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 96638 76074
rect 96690 76022 96742 76074
rect 96794 76022 96846 76074
rect 96898 76022 127358 76074
rect 127410 76022 127462 76074
rect 127514 76022 127566 76074
rect 127618 76022 158078 76074
rect 158130 76022 158182 76074
rect 158234 76022 158286 76074
rect 158338 76022 178640 76074
rect 1344 75988 178640 76022
rect 1344 75290 178640 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 81278 75290
rect 81330 75238 81382 75290
rect 81434 75238 81486 75290
rect 81538 75238 111998 75290
rect 112050 75238 112102 75290
rect 112154 75238 112206 75290
rect 112258 75238 142718 75290
rect 142770 75238 142822 75290
rect 142874 75238 142926 75290
rect 142978 75238 173438 75290
rect 173490 75238 173542 75290
rect 173594 75238 173646 75290
rect 173698 75238 178640 75290
rect 1344 75204 178640 75238
rect 1344 74506 178640 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 96638 74506
rect 96690 74454 96742 74506
rect 96794 74454 96846 74506
rect 96898 74454 127358 74506
rect 127410 74454 127462 74506
rect 127514 74454 127566 74506
rect 127618 74454 158078 74506
rect 158130 74454 158182 74506
rect 158234 74454 158286 74506
rect 158338 74454 178640 74506
rect 1344 74420 178640 74454
rect 1344 73722 178640 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 81278 73722
rect 81330 73670 81382 73722
rect 81434 73670 81486 73722
rect 81538 73670 111998 73722
rect 112050 73670 112102 73722
rect 112154 73670 112206 73722
rect 112258 73670 142718 73722
rect 142770 73670 142822 73722
rect 142874 73670 142926 73722
rect 142978 73670 173438 73722
rect 173490 73670 173542 73722
rect 173594 73670 173646 73722
rect 173698 73670 178640 73722
rect 1344 73636 178640 73670
rect 1344 72938 178640 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 96638 72938
rect 96690 72886 96742 72938
rect 96794 72886 96846 72938
rect 96898 72886 127358 72938
rect 127410 72886 127462 72938
rect 127514 72886 127566 72938
rect 127618 72886 158078 72938
rect 158130 72886 158182 72938
rect 158234 72886 158286 72938
rect 158338 72886 178640 72938
rect 1344 72852 178640 72886
rect 1344 72154 178640 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 81278 72154
rect 81330 72102 81382 72154
rect 81434 72102 81486 72154
rect 81538 72102 111998 72154
rect 112050 72102 112102 72154
rect 112154 72102 112206 72154
rect 112258 72102 142718 72154
rect 142770 72102 142822 72154
rect 142874 72102 142926 72154
rect 142978 72102 173438 72154
rect 173490 72102 173542 72154
rect 173594 72102 173646 72154
rect 173698 72102 178640 72154
rect 1344 72068 178640 72102
rect 1344 71370 178640 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 96638 71370
rect 96690 71318 96742 71370
rect 96794 71318 96846 71370
rect 96898 71318 127358 71370
rect 127410 71318 127462 71370
rect 127514 71318 127566 71370
rect 127618 71318 158078 71370
rect 158130 71318 158182 71370
rect 158234 71318 158286 71370
rect 158338 71318 178640 71370
rect 1344 71284 178640 71318
rect 1344 70586 178640 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 81278 70586
rect 81330 70534 81382 70586
rect 81434 70534 81486 70586
rect 81538 70534 111998 70586
rect 112050 70534 112102 70586
rect 112154 70534 112206 70586
rect 112258 70534 142718 70586
rect 142770 70534 142822 70586
rect 142874 70534 142926 70586
rect 142978 70534 173438 70586
rect 173490 70534 173542 70586
rect 173594 70534 173646 70586
rect 173698 70534 178640 70586
rect 1344 70500 178640 70534
rect 1344 69802 178640 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 96638 69802
rect 96690 69750 96742 69802
rect 96794 69750 96846 69802
rect 96898 69750 127358 69802
rect 127410 69750 127462 69802
rect 127514 69750 127566 69802
rect 127618 69750 158078 69802
rect 158130 69750 158182 69802
rect 158234 69750 158286 69802
rect 158338 69750 178640 69802
rect 1344 69716 178640 69750
rect 1344 69018 178640 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 81278 69018
rect 81330 68966 81382 69018
rect 81434 68966 81486 69018
rect 81538 68966 111998 69018
rect 112050 68966 112102 69018
rect 112154 68966 112206 69018
rect 112258 68966 142718 69018
rect 142770 68966 142822 69018
rect 142874 68966 142926 69018
rect 142978 68966 173438 69018
rect 173490 68966 173542 69018
rect 173594 68966 173646 69018
rect 173698 68966 178640 69018
rect 1344 68932 178640 68966
rect 1344 68234 178640 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 96638 68234
rect 96690 68182 96742 68234
rect 96794 68182 96846 68234
rect 96898 68182 127358 68234
rect 127410 68182 127462 68234
rect 127514 68182 127566 68234
rect 127618 68182 158078 68234
rect 158130 68182 158182 68234
rect 158234 68182 158286 68234
rect 158338 68182 178640 68234
rect 1344 68148 178640 68182
rect 1344 67450 178640 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 81278 67450
rect 81330 67398 81382 67450
rect 81434 67398 81486 67450
rect 81538 67398 111998 67450
rect 112050 67398 112102 67450
rect 112154 67398 112206 67450
rect 112258 67398 142718 67450
rect 142770 67398 142822 67450
rect 142874 67398 142926 67450
rect 142978 67398 173438 67450
rect 173490 67398 173542 67450
rect 173594 67398 173646 67450
rect 173698 67398 178640 67450
rect 1344 67364 178640 67398
rect 1344 66666 178640 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 96638 66666
rect 96690 66614 96742 66666
rect 96794 66614 96846 66666
rect 96898 66614 127358 66666
rect 127410 66614 127462 66666
rect 127514 66614 127566 66666
rect 127618 66614 158078 66666
rect 158130 66614 158182 66666
rect 158234 66614 158286 66666
rect 158338 66614 178640 66666
rect 1344 66580 178640 66614
rect 1344 65882 178640 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 81278 65882
rect 81330 65830 81382 65882
rect 81434 65830 81486 65882
rect 81538 65830 111998 65882
rect 112050 65830 112102 65882
rect 112154 65830 112206 65882
rect 112258 65830 142718 65882
rect 142770 65830 142822 65882
rect 142874 65830 142926 65882
rect 142978 65830 173438 65882
rect 173490 65830 173542 65882
rect 173594 65830 173646 65882
rect 173698 65830 178640 65882
rect 1344 65796 178640 65830
rect 1344 65098 178640 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 96638 65098
rect 96690 65046 96742 65098
rect 96794 65046 96846 65098
rect 96898 65046 127358 65098
rect 127410 65046 127462 65098
rect 127514 65046 127566 65098
rect 127618 65046 158078 65098
rect 158130 65046 158182 65098
rect 158234 65046 158286 65098
rect 158338 65046 178640 65098
rect 1344 65012 178640 65046
rect 1344 64314 178640 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 81278 64314
rect 81330 64262 81382 64314
rect 81434 64262 81486 64314
rect 81538 64262 111998 64314
rect 112050 64262 112102 64314
rect 112154 64262 112206 64314
rect 112258 64262 142718 64314
rect 142770 64262 142822 64314
rect 142874 64262 142926 64314
rect 142978 64262 173438 64314
rect 173490 64262 173542 64314
rect 173594 64262 173646 64314
rect 173698 64262 178640 64314
rect 1344 64228 178640 64262
rect 1344 63530 178640 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 96638 63530
rect 96690 63478 96742 63530
rect 96794 63478 96846 63530
rect 96898 63478 127358 63530
rect 127410 63478 127462 63530
rect 127514 63478 127566 63530
rect 127618 63478 158078 63530
rect 158130 63478 158182 63530
rect 158234 63478 158286 63530
rect 158338 63478 178640 63530
rect 1344 63444 178640 63478
rect 1344 62746 178640 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 81278 62746
rect 81330 62694 81382 62746
rect 81434 62694 81486 62746
rect 81538 62694 111998 62746
rect 112050 62694 112102 62746
rect 112154 62694 112206 62746
rect 112258 62694 142718 62746
rect 142770 62694 142822 62746
rect 142874 62694 142926 62746
rect 142978 62694 173438 62746
rect 173490 62694 173542 62746
rect 173594 62694 173646 62746
rect 173698 62694 178640 62746
rect 1344 62660 178640 62694
rect 1344 61962 178640 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 96638 61962
rect 96690 61910 96742 61962
rect 96794 61910 96846 61962
rect 96898 61910 127358 61962
rect 127410 61910 127462 61962
rect 127514 61910 127566 61962
rect 127618 61910 158078 61962
rect 158130 61910 158182 61962
rect 158234 61910 158286 61962
rect 158338 61910 178640 61962
rect 1344 61876 178640 61910
rect 1344 61178 178640 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 81278 61178
rect 81330 61126 81382 61178
rect 81434 61126 81486 61178
rect 81538 61126 111998 61178
rect 112050 61126 112102 61178
rect 112154 61126 112206 61178
rect 112258 61126 142718 61178
rect 142770 61126 142822 61178
rect 142874 61126 142926 61178
rect 142978 61126 173438 61178
rect 173490 61126 173542 61178
rect 173594 61126 173646 61178
rect 173698 61126 178640 61178
rect 1344 61092 178640 61126
rect 1344 60394 178640 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 96638 60394
rect 96690 60342 96742 60394
rect 96794 60342 96846 60394
rect 96898 60342 127358 60394
rect 127410 60342 127462 60394
rect 127514 60342 127566 60394
rect 127618 60342 158078 60394
rect 158130 60342 158182 60394
rect 158234 60342 158286 60394
rect 158338 60342 178640 60394
rect 1344 60308 178640 60342
rect 1344 59610 178640 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 81278 59610
rect 81330 59558 81382 59610
rect 81434 59558 81486 59610
rect 81538 59558 111998 59610
rect 112050 59558 112102 59610
rect 112154 59558 112206 59610
rect 112258 59558 142718 59610
rect 142770 59558 142822 59610
rect 142874 59558 142926 59610
rect 142978 59558 173438 59610
rect 173490 59558 173542 59610
rect 173594 59558 173646 59610
rect 173698 59558 178640 59610
rect 1344 59524 178640 59558
rect 1344 58826 178640 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 96638 58826
rect 96690 58774 96742 58826
rect 96794 58774 96846 58826
rect 96898 58774 127358 58826
rect 127410 58774 127462 58826
rect 127514 58774 127566 58826
rect 127618 58774 158078 58826
rect 158130 58774 158182 58826
rect 158234 58774 158286 58826
rect 158338 58774 178640 58826
rect 1344 58740 178640 58774
rect 1344 58042 178640 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 81278 58042
rect 81330 57990 81382 58042
rect 81434 57990 81486 58042
rect 81538 57990 111998 58042
rect 112050 57990 112102 58042
rect 112154 57990 112206 58042
rect 112258 57990 142718 58042
rect 142770 57990 142822 58042
rect 142874 57990 142926 58042
rect 142978 57990 173438 58042
rect 173490 57990 173542 58042
rect 173594 57990 173646 58042
rect 173698 57990 178640 58042
rect 1344 57956 178640 57990
rect 1344 57258 178640 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 96638 57258
rect 96690 57206 96742 57258
rect 96794 57206 96846 57258
rect 96898 57206 127358 57258
rect 127410 57206 127462 57258
rect 127514 57206 127566 57258
rect 127618 57206 158078 57258
rect 158130 57206 158182 57258
rect 158234 57206 158286 57258
rect 158338 57206 178640 57258
rect 1344 57172 178640 57206
rect 1344 56474 178640 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 81278 56474
rect 81330 56422 81382 56474
rect 81434 56422 81486 56474
rect 81538 56422 111998 56474
rect 112050 56422 112102 56474
rect 112154 56422 112206 56474
rect 112258 56422 142718 56474
rect 142770 56422 142822 56474
rect 142874 56422 142926 56474
rect 142978 56422 173438 56474
rect 173490 56422 173542 56474
rect 173594 56422 173646 56474
rect 173698 56422 178640 56474
rect 1344 56388 178640 56422
rect 1344 55690 178640 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 96638 55690
rect 96690 55638 96742 55690
rect 96794 55638 96846 55690
rect 96898 55638 127358 55690
rect 127410 55638 127462 55690
rect 127514 55638 127566 55690
rect 127618 55638 158078 55690
rect 158130 55638 158182 55690
rect 158234 55638 158286 55690
rect 158338 55638 178640 55690
rect 1344 55604 178640 55638
rect 1344 54906 178640 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 81278 54906
rect 81330 54854 81382 54906
rect 81434 54854 81486 54906
rect 81538 54854 111998 54906
rect 112050 54854 112102 54906
rect 112154 54854 112206 54906
rect 112258 54854 142718 54906
rect 142770 54854 142822 54906
rect 142874 54854 142926 54906
rect 142978 54854 173438 54906
rect 173490 54854 173542 54906
rect 173594 54854 173646 54906
rect 173698 54854 178640 54906
rect 1344 54820 178640 54854
rect 1344 54122 178640 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 96638 54122
rect 96690 54070 96742 54122
rect 96794 54070 96846 54122
rect 96898 54070 127358 54122
rect 127410 54070 127462 54122
rect 127514 54070 127566 54122
rect 127618 54070 158078 54122
rect 158130 54070 158182 54122
rect 158234 54070 158286 54122
rect 158338 54070 178640 54122
rect 1344 54036 178640 54070
rect 1344 53338 178640 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 81278 53338
rect 81330 53286 81382 53338
rect 81434 53286 81486 53338
rect 81538 53286 111998 53338
rect 112050 53286 112102 53338
rect 112154 53286 112206 53338
rect 112258 53286 142718 53338
rect 142770 53286 142822 53338
rect 142874 53286 142926 53338
rect 142978 53286 173438 53338
rect 173490 53286 173542 53338
rect 173594 53286 173646 53338
rect 173698 53286 178640 53338
rect 1344 53252 178640 53286
rect 1344 52554 178640 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 96638 52554
rect 96690 52502 96742 52554
rect 96794 52502 96846 52554
rect 96898 52502 127358 52554
rect 127410 52502 127462 52554
rect 127514 52502 127566 52554
rect 127618 52502 158078 52554
rect 158130 52502 158182 52554
rect 158234 52502 158286 52554
rect 158338 52502 178640 52554
rect 1344 52468 178640 52502
rect 1344 51770 178640 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 81278 51770
rect 81330 51718 81382 51770
rect 81434 51718 81486 51770
rect 81538 51718 111998 51770
rect 112050 51718 112102 51770
rect 112154 51718 112206 51770
rect 112258 51718 142718 51770
rect 142770 51718 142822 51770
rect 142874 51718 142926 51770
rect 142978 51718 173438 51770
rect 173490 51718 173542 51770
rect 173594 51718 173646 51770
rect 173698 51718 178640 51770
rect 1344 51684 178640 51718
rect 1344 50986 178640 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 96638 50986
rect 96690 50934 96742 50986
rect 96794 50934 96846 50986
rect 96898 50934 127358 50986
rect 127410 50934 127462 50986
rect 127514 50934 127566 50986
rect 127618 50934 158078 50986
rect 158130 50934 158182 50986
rect 158234 50934 158286 50986
rect 158338 50934 178640 50986
rect 1344 50900 178640 50934
rect 1344 50202 178640 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 81278 50202
rect 81330 50150 81382 50202
rect 81434 50150 81486 50202
rect 81538 50150 111998 50202
rect 112050 50150 112102 50202
rect 112154 50150 112206 50202
rect 112258 50150 142718 50202
rect 142770 50150 142822 50202
rect 142874 50150 142926 50202
rect 142978 50150 173438 50202
rect 173490 50150 173542 50202
rect 173594 50150 173646 50202
rect 173698 50150 178640 50202
rect 1344 50116 178640 50150
rect 1344 49418 178640 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 96638 49418
rect 96690 49366 96742 49418
rect 96794 49366 96846 49418
rect 96898 49366 127358 49418
rect 127410 49366 127462 49418
rect 127514 49366 127566 49418
rect 127618 49366 158078 49418
rect 158130 49366 158182 49418
rect 158234 49366 158286 49418
rect 158338 49366 178640 49418
rect 1344 49332 178640 49366
rect 1344 48634 178640 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 81278 48634
rect 81330 48582 81382 48634
rect 81434 48582 81486 48634
rect 81538 48582 111998 48634
rect 112050 48582 112102 48634
rect 112154 48582 112206 48634
rect 112258 48582 142718 48634
rect 142770 48582 142822 48634
rect 142874 48582 142926 48634
rect 142978 48582 173438 48634
rect 173490 48582 173542 48634
rect 173594 48582 173646 48634
rect 173698 48582 178640 48634
rect 1344 48548 178640 48582
rect 1344 47850 178640 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 96638 47850
rect 96690 47798 96742 47850
rect 96794 47798 96846 47850
rect 96898 47798 127358 47850
rect 127410 47798 127462 47850
rect 127514 47798 127566 47850
rect 127618 47798 158078 47850
rect 158130 47798 158182 47850
rect 158234 47798 158286 47850
rect 158338 47798 178640 47850
rect 1344 47764 178640 47798
rect 1344 47066 178640 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 81278 47066
rect 81330 47014 81382 47066
rect 81434 47014 81486 47066
rect 81538 47014 111998 47066
rect 112050 47014 112102 47066
rect 112154 47014 112206 47066
rect 112258 47014 142718 47066
rect 142770 47014 142822 47066
rect 142874 47014 142926 47066
rect 142978 47014 173438 47066
rect 173490 47014 173542 47066
rect 173594 47014 173646 47066
rect 173698 47014 178640 47066
rect 1344 46980 178640 47014
rect 1344 46282 178640 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 96638 46282
rect 96690 46230 96742 46282
rect 96794 46230 96846 46282
rect 96898 46230 127358 46282
rect 127410 46230 127462 46282
rect 127514 46230 127566 46282
rect 127618 46230 158078 46282
rect 158130 46230 158182 46282
rect 158234 46230 158286 46282
rect 158338 46230 178640 46282
rect 1344 46196 178640 46230
rect 1344 45498 178640 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 81278 45498
rect 81330 45446 81382 45498
rect 81434 45446 81486 45498
rect 81538 45446 111998 45498
rect 112050 45446 112102 45498
rect 112154 45446 112206 45498
rect 112258 45446 142718 45498
rect 142770 45446 142822 45498
rect 142874 45446 142926 45498
rect 142978 45446 173438 45498
rect 173490 45446 173542 45498
rect 173594 45446 173646 45498
rect 173698 45446 178640 45498
rect 1344 45412 178640 45446
rect 1344 44714 178640 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 96638 44714
rect 96690 44662 96742 44714
rect 96794 44662 96846 44714
rect 96898 44662 127358 44714
rect 127410 44662 127462 44714
rect 127514 44662 127566 44714
rect 127618 44662 158078 44714
rect 158130 44662 158182 44714
rect 158234 44662 158286 44714
rect 158338 44662 178640 44714
rect 1344 44628 178640 44662
rect 1344 43930 178640 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 81278 43930
rect 81330 43878 81382 43930
rect 81434 43878 81486 43930
rect 81538 43878 111998 43930
rect 112050 43878 112102 43930
rect 112154 43878 112206 43930
rect 112258 43878 142718 43930
rect 142770 43878 142822 43930
rect 142874 43878 142926 43930
rect 142978 43878 173438 43930
rect 173490 43878 173542 43930
rect 173594 43878 173646 43930
rect 173698 43878 178640 43930
rect 1344 43844 178640 43878
rect 1344 43146 178640 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 96638 43146
rect 96690 43094 96742 43146
rect 96794 43094 96846 43146
rect 96898 43094 127358 43146
rect 127410 43094 127462 43146
rect 127514 43094 127566 43146
rect 127618 43094 158078 43146
rect 158130 43094 158182 43146
rect 158234 43094 158286 43146
rect 158338 43094 178640 43146
rect 1344 43060 178640 43094
rect 1344 42362 178640 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 81278 42362
rect 81330 42310 81382 42362
rect 81434 42310 81486 42362
rect 81538 42310 111998 42362
rect 112050 42310 112102 42362
rect 112154 42310 112206 42362
rect 112258 42310 142718 42362
rect 142770 42310 142822 42362
rect 142874 42310 142926 42362
rect 142978 42310 173438 42362
rect 173490 42310 173542 42362
rect 173594 42310 173646 42362
rect 173698 42310 178640 42362
rect 1344 42276 178640 42310
rect 1344 41578 178640 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 96638 41578
rect 96690 41526 96742 41578
rect 96794 41526 96846 41578
rect 96898 41526 127358 41578
rect 127410 41526 127462 41578
rect 127514 41526 127566 41578
rect 127618 41526 158078 41578
rect 158130 41526 158182 41578
rect 158234 41526 158286 41578
rect 158338 41526 178640 41578
rect 1344 41492 178640 41526
rect 1344 40794 178640 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 81278 40794
rect 81330 40742 81382 40794
rect 81434 40742 81486 40794
rect 81538 40742 111998 40794
rect 112050 40742 112102 40794
rect 112154 40742 112206 40794
rect 112258 40742 142718 40794
rect 142770 40742 142822 40794
rect 142874 40742 142926 40794
rect 142978 40742 173438 40794
rect 173490 40742 173542 40794
rect 173594 40742 173646 40794
rect 173698 40742 178640 40794
rect 1344 40708 178640 40742
rect 1344 40010 178640 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 96638 40010
rect 96690 39958 96742 40010
rect 96794 39958 96846 40010
rect 96898 39958 127358 40010
rect 127410 39958 127462 40010
rect 127514 39958 127566 40010
rect 127618 39958 158078 40010
rect 158130 39958 158182 40010
rect 158234 39958 158286 40010
rect 158338 39958 178640 40010
rect 1344 39924 178640 39958
rect 1344 39226 178640 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 81278 39226
rect 81330 39174 81382 39226
rect 81434 39174 81486 39226
rect 81538 39174 111998 39226
rect 112050 39174 112102 39226
rect 112154 39174 112206 39226
rect 112258 39174 142718 39226
rect 142770 39174 142822 39226
rect 142874 39174 142926 39226
rect 142978 39174 173438 39226
rect 173490 39174 173542 39226
rect 173594 39174 173646 39226
rect 173698 39174 178640 39226
rect 1344 39140 178640 39174
rect 1344 38442 178640 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 96638 38442
rect 96690 38390 96742 38442
rect 96794 38390 96846 38442
rect 96898 38390 127358 38442
rect 127410 38390 127462 38442
rect 127514 38390 127566 38442
rect 127618 38390 158078 38442
rect 158130 38390 158182 38442
rect 158234 38390 158286 38442
rect 158338 38390 178640 38442
rect 1344 38356 178640 38390
rect 1344 37658 178640 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 81278 37658
rect 81330 37606 81382 37658
rect 81434 37606 81486 37658
rect 81538 37606 111998 37658
rect 112050 37606 112102 37658
rect 112154 37606 112206 37658
rect 112258 37606 142718 37658
rect 142770 37606 142822 37658
rect 142874 37606 142926 37658
rect 142978 37606 173438 37658
rect 173490 37606 173542 37658
rect 173594 37606 173646 37658
rect 173698 37606 178640 37658
rect 1344 37572 178640 37606
rect 1344 36874 178640 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 96638 36874
rect 96690 36822 96742 36874
rect 96794 36822 96846 36874
rect 96898 36822 127358 36874
rect 127410 36822 127462 36874
rect 127514 36822 127566 36874
rect 127618 36822 158078 36874
rect 158130 36822 158182 36874
rect 158234 36822 158286 36874
rect 158338 36822 178640 36874
rect 1344 36788 178640 36822
rect 1344 36090 178640 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 81278 36090
rect 81330 36038 81382 36090
rect 81434 36038 81486 36090
rect 81538 36038 111998 36090
rect 112050 36038 112102 36090
rect 112154 36038 112206 36090
rect 112258 36038 142718 36090
rect 142770 36038 142822 36090
rect 142874 36038 142926 36090
rect 142978 36038 173438 36090
rect 173490 36038 173542 36090
rect 173594 36038 173646 36090
rect 173698 36038 178640 36090
rect 1344 36004 178640 36038
rect 1344 35306 178640 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 96638 35306
rect 96690 35254 96742 35306
rect 96794 35254 96846 35306
rect 96898 35254 127358 35306
rect 127410 35254 127462 35306
rect 127514 35254 127566 35306
rect 127618 35254 158078 35306
rect 158130 35254 158182 35306
rect 158234 35254 158286 35306
rect 158338 35254 178640 35306
rect 1344 35220 178640 35254
rect 1344 34522 178640 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 81278 34522
rect 81330 34470 81382 34522
rect 81434 34470 81486 34522
rect 81538 34470 111998 34522
rect 112050 34470 112102 34522
rect 112154 34470 112206 34522
rect 112258 34470 142718 34522
rect 142770 34470 142822 34522
rect 142874 34470 142926 34522
rect 142978 34470 173438 34522
rect 173490 34470 173542 34522
rect 173594 34470 173646 34522
rect 173698 34470 178640 34522
rect 1344 34436 178640 34470
rect 1344 33738 178640 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 96638 33738
rect 96690 33686 96742 33738
rect 96794 33686 96846 33738
rect 96898 33686 127358 33738
rect 127410 33686 127462 33738
rect 127514 33686 127566 33738
rect 127618 33686 158078 33738
rect 158130 33686 158182 33738
rect 158234 33686 158286 33738
rect 158338 33686 178640 33738
rect 1344 33652 178640 33686
rect 1344 32954 178640 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 81278 32954
rect 81330 32902 81382 32954
rect 81434 32902 81486 32954
rect 81538 32902 111998 32954
rect 112050 32902 112102 32954
rect 112154 32902 112206 32954
rect 112258 32902 142718 32954
rect 142770 32902 142822 32954
rect 142874 32902 142926 32954
rect 142978 32902 173438 32954
rect 173490 32902 173542 32954
rect 173594 32902 173646 32954
rect 173698 32902 178640 32954
rect 1344 32868 178640 32902
rect 1344 32170 178640 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 96638 32170
rect 96690 32118 96742 32170
rect 96794 32118 96846 32170
rect 96898 32118 127358 32170
rect 127410 32118 127462 32170
rect 127514 32118 127566 32170
rect 127618 32118 158078 32170
rect 158130 32118 158182 32170
rect 158234 32118 158286 32170
rect 158338 32118 178640 32170
rect 1344 32084 178640 32118
rect 1344 31386 178640 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 81278 31386
rect 81330 31334 81382 31386
rect 81434 31334 81486 31386
rect 81538 31334 111998 31386
rect 112050 31334 112102 31386
rect 112154 31334 112206 31386
rect 112258 31334 142718 31386
rect 142770 31334 142822 31386
rect 142874 31334 142926 31386
rect 142978 31334 173438 31386
rect 173490 31334 173542 31386
rect 173594 31334 173646 31386
rect 173698 31334 178640 31386
rect 1344 31300 178640 31334
rect 1344 30602 178640 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 96638 30602
rect 96690 30550 96742 30602
rect 96794 30550 96846 30602
rect 96898 30550 127358 30602
rect 127410 30550 127462 30602
rect 127514 30550 127566 30602
rect 127618 30550 158078 30602
rect 158130 30550 158182 30602
rect 158234 30550 158286 30602
rect 158338 30550 178640 30602
rect 1344 30516 178640 30550
rect 1344 29818 178640 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 81278 29818
rect 81330 29766 81382 29818
rect 81434 29766 81486 29818
rect 81538 29766 111998 29818
rect 112050 29766 112102 29818
rect 112154 29766 112206 29818
rect 112258 29766 142718 29818
rect 142770 29766 142822 29818
rect 142874 29766 142926 29818
rect 142978 29766 173438 29818
rect 173490 29766 173542 29818
rect 173594 29766 173646 29818
rect 173698 29766 178640 29818
rect 1344 29732 178640 29766
rect 1344 29034 178640 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 96638 29034
rect 96690 28982 96742 29034
rect 96794 28982 96846 29034
rect 96898 28982 127358 29034
rect 127410 28982 127462 29034
rect 127514 28982 127566 29034
rect 127618 28982 158078 29034
rect 158130 28982 158182 29034
rect 158234 28982 158286 29034
rect 158338 28982 178640 29034
rect 1344 28948 178640 28982
rect 1344 28250 178640 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 81278 28250
rect 81330 28198 81382 28250
rect 81434 28198 81486 28250
rect 81538 28198 111998 28250
rect 112050 28198 112102 28250
rect 112154 28198 112206 28250
rect 112258 28198 142718 28250
rect 142770 28198 142822 28250
rect 142874 28198 142926 28250
rect 142978 28198 173438 28250
rect 173490 28198 173542 28250
rect 173594 28198 173646 28250
rect 173698 28198 178640 28250
rect 1344 28164 178640 28198
rect 1344 27466 178640 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 96638 27466
rect 96690 27414 96742 27466
rect 96794 27414 96846 27466
rect 96898 27414 127358 27466
rect 127410 27414 127462 27466
rect 127514 27414 127566 27466
rect 127618 27414 158078 27466
rect 158130 27414 158182 27466
rect 158234 27414 158286 27466
rect 158338 27414 178640 27466
rect 1344 27380 178640 27414
rect 1344 26682 178640 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 81278 26682
rect 81330 26630 81382 26682
rect 81434 26630 81486 26682
rect 81538 26630 111998 26682
rect 112050 26630 112102 26682
rect 112154 26630 112206 26682
rect 112258 26630 142718 26682
rect 142770 26630 142822 26682
rect 142874 26630 142926 26682
rect 142978 26630 173438 26682
rect 173490 26630 173542 26682
rect 173594 26630 173646 26682
rect 173698 26630 178640 26682
rect 1344 26596 178640 26630
rect 1344 25898 178640 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 96638 25898
rect 96690 25846 96742 25898
rect 96794 25846 96846 25898
rect 96898 25846 127358 25898
rect 127410 25846 127462 25898
rect 127514 25846 127566 25898
rect 127618 25846 158078 25898
rect 158130 25846 158182 25898
rect 158234 25846 158286 25898
rect 158338 25846 178640 25898
rect 1344 25812 178640 25846
rect 1344 25114 178640 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 81278 25114
rect 81330 25062 81382 25114
rect 81434 25062 81486 25114
rect 81538 25062 111998 25114
rect 112050 25062 112102 25114
rect 112154 25062 112206 25114
rect 112258 25062 142718 25114
rect 142770 25062 142822 25114
rect 142874 25062 142926 25114
rect 142978 25062 173438 25114
rect 173490 25062 173542 25114
rect 173594 25062 173646 25114
rect 173698 25062 178640 25114
rect 1344 25028 178640 25062
rect 1344 24330 178640 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 96638 24330
rect 96690 24278 96742 24330
rect 96794 24278 96846 24330
rect 96898 24278 127358 24330
rect 127410 24278 127462 24330
rect 127514 24278 127566 24330
rect 127618 24278 158078 24330
rect 158130 24278 158182 24330
rect 158234 24278 158286 24330
rect 158338 24278 178640 24330
rect 1344 24244 178640 24278
rect 1344 23546 178640 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 81278 23546
rect 81330 23494 81382 23546
rect 81434 23494 81486 23546
rect 81538 23494 111998 23546
rect 112050 23494 112102 23546
rect 112154 23494 112206 23546
rect 112258 23494 142718 23546
rect 142770 23494 142822 23546
rect 142874 23494 142926 23546
rect 142978 23494 173438 23546
rect 173490 23494 173542 23546
rect 173594 23494 173646 23546
rect 173698 23494 178640 23546
rect 1344 23460 178640 23494
rect 1344 22762 178640 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 96638 22762
rect 96690 22710 96742 22762
rect 96794 22710 96846 22762
rect 96898 22710 127358 22762
rect 127410 22710 127462 22762
rect 127514 22710 127566 22762
rect 127618 22710 158078 22762
rect 158130 22710 158182 22762
rect 158234 22710 158286 22762
rect 158338 22710 178640 22762
rect 1344 22676 178640 22710
rect 1344 21978 178640 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 81278 21978
rect 81330 21926 81382 21978
rect 81434 21926 81486 21978
rect 81538 21926 111998 21978
rect 112050 21926 112102 21978
rect 112154 21926 112206 21978
rect 112258 21926 142718 21978
rect 142770 21926 142822 21978
rect 142874 21926 142926 21978
rect 142978 21926 173438 21978
rect 173490 21926 173542 21978
rect 173594 21926 173646 21978
rect 173698 21926 178640 21978
rect 1344 21892 178640 21926
rect 1344 21194 178640 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 96638 21194
rect 96690 21142 96742 21194
rect 96794 21142 96846 21194
rect 96898 21142 127358 21194
rect 127410 21142 127462 21194
rect 127514 21142 127566 21194
rect 127618 21142 158078 21194
rect 158130 21142 158182 21194
rect 158234 21142 158286 21194
rect 158338 21142 178640 21194
rect 1344 21108 178640 21142
rect 1344 20410 178640 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 81278 20410
rect 81330 20358 81382 20410
rect 81434 20358 81486 20410
rect 81538 20358 111998 20410
rect 112050 20358 112102 20410
rect 112154 20358 112206 20410
rect 112258 20358 142718 20410
rect 142770 20358 142822 20410
rect 142874 20358 142926 20410
rect 142978 20358 173438 20410
rect 173490 20358 173542 20410
rect 173594 20358 173646 20410
rect 173698 20358 178640 20410
rect 1344 20324 178640 20358
rect 1344 19626 178640 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 96638 19626
rect 96690 19574 96742 19626
rect 96794 19574 96846 19626
rect 96898 19574 127358 19626
rect 127410 19574 127462 19626
rect 127514 19574 127566 19626
rect 127618 19574 158078 19626
rect 158130 19574 158182 19626
rect 158234 19574 158286 19626
rect 158338 19574 178640 19626
rect 1344 19540 178640 19574
rect 1344 18842 178640 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 81278 18842
rect 81330 18790 81382 18842
rect 81434 18790 81486 18842
rect 81538 18790 111998 18842
rect 112050 18790 112102 18842
rect 112154 18790 112206 18842
rect 112258 18790 142718 18842
rect 142770 18790 142822 18842
rect 142874 18790 142926 18842
rect 142978 18790 173438 18842
rect 173490 18790 173542 18842
rect 173594 18790 173646 18842
rect 173698 18790 178640 18842
rect 1344 18756 178640 18790
rect 1344 18058 178640 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 96638 18058
rect 96690 18006 96742 18058
rect 96794 18006 96846 18058
rect 96898 18006 127358 18058
rect 127410 18006 127462 18058
rect 127514 18006 127566 18058
rect 127618 18006 158078 18058
rect 158130 18006 158182 18058
rect 158234 18006 158286 18058
rect 158338 18006 178640 18058
rect 1344 17972 178640 18006
rect 1344 17274 178640 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 81278 17274
rect 81330 17222 81382 17274
rect 81434 17222 81486 17274
rect 81538 17222 111998 17274
rect 112050 17222 112102 17274
rect 112154 17222 112206 17274
rect 112258 17222 142718 17274
rect 142770 17222 142822 17274
rect 142874 17222 142926 17274
rect 142978 17222 173438 17274
rect 173490 17222 173542 17274
rect 173594 17222 173646 17274
rect 173698 17222 178640 17274
rect 1344 17188 178640 17222
rect 1344 16490 178640 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 96638 16490
rect 96690 16438 96742 16490
rect 96794 16438 96846 16490
rect 96898 16438 127358 16490
rect 127410 16438 127462 16490
rect 127514 16438 127566 16490
rect 127618 16438 158078 16490
rect 158130 16438 158182 16490
rect 158234 16438 158286 16490
rect 158338 16438 178640 16490
rect 1344 16404 178640 16438
rect 1344 15706 178640 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 81278 15706
rect 81330 15654 81382 15706
rect 81434 15654 81486 15706
rect 81538 15654 111998 15706
rect 112050 15654 112102 15706
rect 112154 15654 112206 15706
rect 112258 15654 142718 15706
rect 142770 15654 142822 15706
rect 142874 15654 142926 15706
rect 142978 15654 173438 15706
rect 173490 15654 173542 15706
rect 173594 15654 173646 15706
rect 173698 15654 178640 15706
rect 1344 15620 178640 15654
rect 1344 14922 178640 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 96638 14922
rect 96690 14870 96742 14922
rect 96794 14870 96846 14922
rect 96898 14870 127358 14922
rect 127410 14870 127462 14922
rect 127514 14870 127566 14922
rect 127618 14870 158078 14922
rect 158130 14870 158182 14922
rect 158234 14870 158286 14922
rect 158338 14870 178640 14922
rect 1344 14836 178640 14870
rect 1344 14138 178640 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 81278 14138
rect 81330 14086 81382 14138
rect 81434 14086 81486 14138
rect 81538 14086 111998 14138
rect 112050 14086 112102 14138
rect 112154 14086 112206 14138
rect 112258 14086 142718 14138
rect 142770 14086 142822 14138
rect 142874 14086 142926 14138
rect 142978 14086 173438 14138
rect 173490 14086 173542 14138
rect 173594 14086 173646 14138
rect 173698 14086 178640 14138
rect 1344 14052 178640 14086
rect 69134 13634 69186 13646
rect 69134 13570 69186 13582
rect 69582 13634 69634 13646
rect 69582 13570 69634 13582
rect 70030 13634 70082 13646
rect 70030 13570 70082 13582
rect 70590 13634 70642 13646
rect 70590 13570 70642 13582
rect 71038 13634 71090 13646
rect 71038 13570 71090 13582
rect 72718 13634 72770 13646
rect 72718 13570 72770 13582
rect 74958 13634 75010 13646
rect 74958 13570 75010 13582
rect 75406 13634 75458 13646
rect 75406 13570 75458 13582
rect 75854 13634 75906 13646
rect 75854 13570 75906 13582
rect 77086 13634 77138 13646
rect 77086 13570 77138 13582
rect 78206 13634 78258 13646
rect 78206 13570 78258 13582
rect 79102 13634 79154 13646
rect 79102 13570 79154 13582
rect 79774 13634 79826 13646
rect 79774 13570 79826 13582
rect 80670 13634 80722 13646
rect 80670 13570 80722 13582
rect 1344 13354 178640 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 96638 13354
rect 96690 13302 96742 13354
rect 96794 13302 96846 13354
rect 96898 13302 127358 13354
rect 127410 13302 127462 13354
rect 127514 13302 127566 13354
rect 127618 13302 158078 13354
rect 158130 13302 158182 13354
rect 158234 13302 158286 13354
rect 158338 13302 178640 13354
rect 1344 13268 178640 13302
rect 75730 13134 75742 13186
rect 75794 13183 75806 13186
rect 76402 13183 76414 13186
rect 75794 13137 76414 13183
rect 75794 13134 75806 13137
rect 76402 13134 76414 13137
rect 76466 13134 76478 13186
rect 79202 13134 79214 13186
rect 79266 13183 79278 13186
rect 79538 13183 79550 13186
rect 79266 13137 79550 13183
rect 79266 13134 79278 13137
rect 79538 13134 79550 13137
rect 79602 13183 79614 13186
rect 79762 13183 79774 13186
rect 79602 13137 79774 13183
rect 79602 13134 79614 13137
rect 79762 13134 79774 13137
rect 79826 13134 79838 13186
rect 68238 13074 68290 13086
rect 68238 13010 68290 13022
rect 69694 13074 69746 13086
rect 69694 13010 69746 13022
rect 70142 13074 70194 13086
rect 70142 13010 70194 13022
rect 71262 13074 71314 13086
rect 71262 13010 71314 13022
rect 72270 13074 72322 13086
rect 72270 13010 72322 13022
rect 73502 13074 73554 13086
rect 73502 13010 73554 13022
rect 75742 13074 75794 13086
rect 75742 13010 75794 13022
rect 83022 13074 83074 13086
rect 104066 13022 104078 13074
rect 104130 13022 104142 13074
rect 83022 13010 83074 13022
rect 76638 12962 76690 12974
rect 101154 12910 101166 12962
rect 101218 12910 101230 12962
rect 76638 12898 76690 12910
rect 79662 12850 79714 12862
rect 101938 12798 101950 12850
rect 102002 12798 102014 12850
rect 79662 12786 79714 12798
rect 67342 12738 67394 12750
rect 67342 12674 67394 12686
rect 68686 12738 68738 12750
rect 68686 12674 68738 12686
rect 70814 12738 70866 12750
rect 70814 12674 70866 12686
rect 71710 12738 71762 12750
rect 71710 12674 71762 12686
rect 72718 12738 72770 12750
rect 72718 12674 72770 12686
rect 73166 12738 73218 12750
rect 73166 12674 73218 12686
rect 74174 12738 74226 12750
rect 74174 12674 74226 12686
rect 74734 12738 74786 12750
rect 74734 12674 74786 12686
rect 75182 12738 75234 12750
rect 75182 12674 75234 12686
rect 76190 12738 76242 12750
rect 76190 12674 76242 12686
rect 77198 12738 77250 12750
rect 77198 12674 77250 12686
rect 77758 12738 77810 12750
rect 77758 12674 77810 12686
rect 78542 12738 78594 12750
rect 78542 12674 78594 12686
rect 79102 12738 79154 12750
rect 79102 12674 79154 12686
rect 79998 12738 80050 12750
rect 79998 12674 80050 12686
rect 80894 12738 80946 12750
rect 80894 12674 80946 12686
rect 81454 12738 81506 12750
rect 81454 12674 81506 12686
rect 82686 12738 82738 12750
rect 82686 12674 82738 12686
rect 100382 12738 100434 12750
rect 100382 12674 100434 12686
rect 1344 12570 178640 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 81278 12570
rect 81330 12518 81382 12570
rect 81434 12518 81486 12570
rect 81538 12518 111998 12570
rect 112050 12518 112102 12570
rect 112154 12518 112206 12570
rect 112258 12518 142718 12570
rect 142770 12518 142822 12570
rect 142874 12518 142926 12570
rect 142978 12518 173438 12570
rect 173490 12518 173542 12570
rect 173594 12518 173646 12570
rect 173698 12518 178640 12570
rect 1344 12484 178640 12518
rect 52782 12402 52834 12414
rect 52782 12338 52834 12350
rect 57934 12402 57986 12414
rect 57934 12338 57986 12350
rect 64206 12402 64258 12414
rect 64206 12338 64258 12350
rect 70254 12402 70306 12414
rect 70254 12338 70306 12350
rect 76078 12402 76130 12414
rect 76078 12338 76130 12350
rect 76526 12402 76578 12414
rect 76526 12338 76578 12350
rect 77086 12402 77138 12414
rect 77086 12338 77138 12350
rect 77422 12402 77474 12414
rect 77422 12338 77474 12350
rect 77982 12402 78034 12414
rect 77982 12338 78034 12350
rect 79214 12402 79266 12414
rect 79214 12338 79266 12350
rect 80558 12402 80610 12414
rect 80558 12338 80610 12350
rect 81678 12402 81730 12414
rect 81678 12338 81730 12350
rect 82574 12402 82626 12414
rect 82574 12338 82626 12350
rect 85934 12402 85986 12414
rect 85934 12338 85986 12350
rect 57374 12290 57426 12302
rect 57374 12226 57426 12238
rect 59614 12290 59666 12302
rect 63758 12290 63810 12302
rect 60834 12238 60846 12290
rect 60898 12238 60910 12290
rect 61170 12238 61182 12290
rect 61234 12238 61246 12290
rect 59614 12226 59666 12238
rect 63758 12226 63810 12238
rect 73614 12290 73666 12302
rect 73614 12226 73666 12238
rect 91086 12290 91138 12302
rect 91086 12226 91138 12238
rect 91198 12178 91250 12190
rect 98802 12126 98814 12178
rect 98866 12126 98878 12178
rect 105186 12126 105198 12178
rect 105250 12126 105262 12178
rect 108658 12126 108670 12178
rect 108722 12126 108734 12178
rect 91198 12114 91250 12126
rect 55134 12066 55186 12078
rect 55134 12002 55186 12014
rect 58382 12066 58434 12078
rect 58382 12002 58434 12014
rect 59166 12066 59218 12078
rect 59166 12002 59218 12014
rect 61966 12066 62018 12078
rect 61966 12002 62018 12014
rect 64766 12066 64818 12078
rect 64766 12002 64818 12014
rect 65662 12066 65714 12078
rect 65662 12002 65714 12014
rect 66110 12066 66162 12078
rect 66110 12002 66162 12014
rect 66894 12066 66946 12078
rect 66894 12002 66946 12014
rect 67454 12066 67506 12078
rect 67454 12002 67506 12014
rect 68126 12066 68178 12078
rect 68126 12002 68178 12014
rect 68686 12066 68738 12078
rect 68686 12002 68738 12014
rect 69134 12066 69186 12078
rect 69134 12002 69186 12014
rect 69582 12066 69634 12078
rect 69582 12002 69634 12014
rect 70590 12066 70642 12078
rect 70590 12002 70642 12014
rect 71038 12066 71090 12078
rect 71038 12002 71090 12014
rect 71934 12066 71986 12078
rect 71934 12002 71986 12014
rect 72382 12066 72434 12078
rect 72382 12002 72434 12014
rect 74174 12066 74226 12078
rect 74174 12002 74226 12014
rect 74510 12066 74562 12078
rect 74510 12002 74562 12014
rect 74958 12066 75010 12078
rect 74958 12002 75010 12014
rect 75518 12066 75570 12078
rect 75518 12002 75570 12014
rect 78542 12066 78594 12078
rect 78542 12002 78594 12014
rect 79662 12066 79714 12078
rect 79662 12002 79714 12014
rect 80110 12066 80162 12078
rect 80110 12002 80162 12014
rect 81342 12066 81394 12078
rect 81342 12002 81394 12014
rect 82238 12066 82290 12078
rect 82238 12002 82290 12014
rect 83246 12066 83298 12078
rect 83246 12002 83298 12014
rect 83694 12066 83746 12078
rect 83694 12002 83746 12014
rect 84142 12066 84194 12078
rect 84142 12002 84194 12014
rect 84814 12066 84866 12078
rect 84814 12002 84866 12014
rect 90414 12066 90466 12078
rect 90414 12002 90466 12014
rect 98142 12066 98194 12078
rect 101614 12066 101666 12078
rect 99474 12014 99486 12066
rect 99538 12014 99550 12066
rect 98142 12002 98194 12014
rect 101614 12002 101666 12014
rect 104526 12066 104578 12078
rect 112142 12066 112194 12078
rect 105970 12014 105982 12066
rect 106034 12014 106046 12066
rect 108098 12014 108110 12066
rect 108162 12014 108174 12066
rect 109442 12014 109454 12066
rect 109506 12014 109518 12066
rect 111570 12014 111582 12066
rect 111634 12014 111646 12066
rect 104526 12002 104578 12014
rect 112142 12002 112194 12014
rect 60286 11954 60338 11966
rect 57250 11902 57262 11954
rect 57314 11951 57326 11954
rect 58370 11951 58382 11954
rect 57314 11905 58382 11951
rect 57314 11902 57326 11905
rect 58370 11902 58382 11905
rect 58434 11902 58446 11954
rect 60286 11890 60338 11902
rect 60622 11954 60674 11966
rect 91310 11954 91362 11966
rect 68114 11902 68126 11954
rect 68178 11951 68190 11954
rect 68562 11951 68574 11954
rect 68178 11905 68574 11951
rect 68178 11902 68190 11905
rect 68562 11902 68574 11905
rect 68626 11902 68638 11954
rect 60622 11890 60674 11902
rect 91310 11890 91362 11902
rect 1344 11786 178640 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 96638 11786
rect 96690 11734 96742 11786
rect 96794 11734 96846 11786
rect 96898 11734 127358 11786
rect 127410 11734 127462 11786
rect 127514 11734 127566 11786
rect 127618 11734 158078 11786
rect 158130 11734 158182 11786
rect 158234 11734 158286 11786
rect 158338 11734 178640 11786
rect 1344 11700 178640 11734
rect 57138 11566 57150 11618
rect 57202 11615 57214 11618
rect 57922 11615 57934 11618
rect 57202 11569 57934 11615
rect 57202 11566 57214 11569
rect 57922 11566 57934 11569
rect 57986 11566 57998 11618
rect 99810 11566 99822 11618
rect 99874 11615 99886 11618
rect 100594 11615 100606 11618
rect 99874 11569 100606 11615
rect 99874 11566 99886 11569
rect 100594 11566 100606 11569
rect 100658 11566 100670 11618
rect 107426 11615 107438 11618
rect 106993 11569 107438 11615
rect 47182 11506 47234 11518
rect 47182 11442 47234 11454
rect 51998 11506 52050 11518
rect 51998 11442 52050 11454
rect 54462 11506 54514 11518
rect 54462 11442 54514 11454
rect 55022 11506 55074 11518
rect 55022 11442 55074 11454
rect 57934 11506 57986 11518
rect 57934 11442 57986 11454
rect 58382 11506 58434 11518
rect 58382 11442 58434 11454
rect 59950 11506 60002 11518
rect 67790 11506 67842 11518
rect 63746 11454 63758 11506
rect 63810 11454 63822 11506
rect 59950 11442 60002 11454
rect 67790 11442 67842 11454
rect 70142 11506 70194 11518
rect 70142 11442 70194 11454
rect 77198 11506 77250 11518
rect 77198 11442 77250 11454
rect 78094 11506 78146 11518
rect 82798 11506 82850 11518
rect 99262 11506 99314 11518
rect 79426 11454 79438 11506
rect 79490 11454 79502 11506
rect 85362 11454 85374 11506
rect 85426 11454 85438 11506
rect 89506 11454 89518 11506
rect 89570 11454 89582 11506
rect 91634 11454 91646 11506
rect 91698 11454 91710 11506
rect 97234 11454 97246 11506
rect 97298 11454 97310 11506
rect 78094 11442 78146 11454
rect 82798 11442 82850 11454
rect 99262 11442 99314 11454
rect 69694 11394 69746 11406
rect 66546 11342 66558 11394
rect 66610 11342 66622 11394
rect 69694 11330 69746 11342
rect 70702 11394 70754 11406
rect 78430 11394 78482 11406
rect 88958 11394 89010 11406
rect 93774 11394 93826 11406
rect 72594 11342 72606 11394
rect 72658 11342 72670 11394
rect 73378 11342 73390 11394
rect 73442 11342 73454 11394
rect 82226 11342 82238 11394
rect 82290 11342 82302 11394
rect 88386 11342 88398 11394
rect 88450 11342 88462 11394
rect 92418 11342 92430 11394
rect 92482 11342 92494 11394
rect 70702 11330 70754 11342
rect 78430 11330 78482 11342
rect 88958 11330 89010 11342
rect 93774 11330 93826 11342
rect 94322 11330 94334 11382
rect 94386 11330 94398 11382
rect 103394 11342 103406 11394
rect 103458 11342 103470 11394
rect 106642 11342 106654 11394
rect 106706 11391 106718 11394
rect 106993 11391 107039 11569
rect 107426 11566 107438 11569
rect 107490 11566 107502 11618
rect 107438 11506 107490 11518
rect 107438 11442 107490 11454
rect 112030 11506 112082 11518
rect 112030 11442 112082 11454
rect 115278 11506 115330 11518
rect 115278 11442 115330 11454
rect 106706 11345 107039 11391
rect 106706 11342 106718 11345
rect 109106 11342 109118 11394
rect 109170 11342 109182 11394
rect 51102 11282 51154 11294
rect 51102 11218 51154 11230
rect 54014 11282 54066 11294
rect 70814 11282 70866 11294
rect 65874 11230 65886 11282
rect 65938 11230 65950 11282
rect 54014 11218 54066 11230
rect 70814 11218 70866 11230
rect 71822 11282 71874 11294
rect 83470 11282 83522 11294
rect 81554 11230 81566 11282
rect 81618 11230 81630 11282
rect 71822 11218 71874 11230
rect 83470 11218 83522 11230
rect 83694 11282 83746 11294
rect 99374 11282 99426 11294
rect 87602 11230 87614 11282
rect 87666 11230 87678 11282
rect 95106 11230 95118 11282
rect 95170 11230 95182 11282
rect 83694 11218 83746 11230
rect 99374 11218 99426 11230
rect 99934 11282 99986 11294
rect 104178 11230 104190 11282
rect 104242 11230 104254 11282
rect 109890 11230 109902 11282
rect 109954 11230 109966 11282
rect 99934 11218 99986 11230
rect 39118 11170 39170 11182
rect 39118 11106 39170 11118
rect 39566 11170 39618 11182
rect 39566 11106 39618 11118
rect 46622 11170 46674 11182
rect 46622 11106 46674 11118
rect 47630 11170 47682 11182
rect 47630 11106 47682 11118
rect 48078 11170 48130 11182
rect 48078 11106 48130 11118
rect 48750 11170 48802 11182
rect 48750 11106 48802 11118
rect 51662 11170 51714 11182
rect 51662 11106 51714 11118
rect 52782 11170 52834 11182
rect 52782 11106 52834 11118
rect 53678 11170 53730 11182
rect 53678 11106 53730 11118
rect 55582 11170 55634 11182
rect 55582 11106 55634 11118
rect 56030 11170 56082 11182
rect 56030 11106 56082 11118
rect 56366 11170 56418 11182
rect 56366 11106 56418 11118
rect 56814 11170 56866 11182
rect 56814 11106 56866 11118
rect 57486 11170 57538 11182
rect 57486 11106 57538 11118
rect 58718 11170 58770 11182
rect 58718 11106 58770 11118
rect 60286 11170 60338 11182
rect 60286 11106 60338 11118
rect 61294 11170 61346 11182
rect 61294 11106 61346 11118
rect 61854 11170 61906 11182
rect 61854 11106 61906 11118
rect 62190 11170 62242 11182
rect 62190 11106 62242 11118
rect 62638 11170 62690 11182
rect 62638 11106 62690 11118
rect 63198 11170 63250 11182
rect 63198 11106 63250 11118
rect 67118 11170 67170 11182
rect 67118 11106 67170 11118
rect 68126 11170 68178 11182
rect 68126 11106 68178 11118
rect 68574 11170 68626 11182
rect 68574 11106 68626 11118
rect 69246 11170 69298 11182
rect 69246 11106 69298 11118
rect 71038 11170 71090 11182
rect 71038 11106 71090 11118
rect 71598 11170 71650 11182
rect 71598 11106 71650 11118
rect 71710 11170 71762 11182
rect 76190 11170 76242 11182
rect 75618 11118 75630 11170
rect 75682 11118 75694 11170
rect 71710 11106 71762 11118
rect 76190 11106 76242 11118
rect 78878 11170 78930 11182
rect 78878 11106 78930 11118
rect 83582 11170 83634 11182
rect 83582 11106 83634 11118
rect 84478 11170 84530 11182
rect 84478 11106 84530 11118
rect 97694 11170 97746 11182
rect 97694 11106 97746 11118
rect 98254 11170 98306 11182
rect 98254 11106 98306 11118
rect 99150 11170 99202 11182
rect 99150 11106 99202 11118
rect 100382 11170 100434 11182
rect 100382 11106 100434 11118
rect 101166 11170 101218 11182
rect 101166 11106 101218 11118
rect 101502 11170 101554 11182
rect 101502 11106 101554 11118
rect 101950 11170 102002 11182
rect 101950 11106 102002 11118
rect 102846 11170 102898 11182
rect 107102 11170 107154 11182
rect 106418 11118 106430 11170
rect 106482 11118 106494 11170
rect 102846 11106 102898 11118
rect 107102 11106 107154 11118
rect 107886 11170 107938 11182
rect 107886 11106 107938 11118
rect 108334 11170 108386 11182
rect 108334 11106 108386 11118
rect 112702 11170 112754 11182
rect 112702 11106 112754 11118
rect 113150 11170 113202 11182
rect 113150 11106 113202 11118
rect 114718 11170 114770 11182
rect 114718 11106 114770 11118
rect 1344 11002 178640 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 81278 11002
rect 81330 10950 81382 11002
rect 81434 10950 81486 11002
rect 81538 10950 111998 11002
rect 112050 10950 112102 11002
rect 112154 10950 112206 11002
rect 112258 10950 142718 11002
rect 142770 10950 142822 11002
rect 142874 10950 142926 11002
rect 142978 10950 173438 11002
rect 173490 10950 173542 11002
rect 173594 10950 173646 11002
rect 173698 10950 178640 11002
rect 1344 10916 178640 10950
rect 39342 10834 39394 10846
rect 39342 10770 39394 10782
rect 46398 10834 46450 10846
rect 46398 10770 46450 10782
rect 48750 10834 48802 10846
rect 48750 10770 48802 10782
rect 56030 10834 56082 10846
rect 56030 10770 56082 10782
rect 63422 10834 63474 10846
rect 63422 10770 63474 10782
rect 65550 10834 65602 10846
rect 65550 10770 65602 10782
rect 74286 10834 74338 10846
rect 74286 10770 74338 10782
rect 75742 10834 75794 10846
rect 82126 10834 82178 10846
rect 76850 10782 76862 10834
rect 76914 10782 76926 10834
rect 75742 10770 75794 10782
rect 82126 10770 82178 10782
rect 86382 10834 86434 10846
rect 86382 10770 86434 10782
rect 96462 10834 96514 10846
rect 96462 10770 96514 10782
rect 100606 10834 100658 10846
rect 100606 10770 100658 10782
rect 101054 10834 101106 10846
rect 101054 10770 101106 10782
rect 101614 10834 101666 10846
rect 101614 10770 101666 10782
rect 104302 10834 104354 10846
rect 104302 10770 104354 10782
rect 105422 10834 105474 10846
rect 105422 10770 105474 10782
rect 106430 10834 106482 10846
rect 106430 10770 106482 10782
rect 108558 10834 108610 10846
rect 108558 10770 108610 10782
rect 115054 10834 115106 10846
rect 115054 10770 115106 10782
rect 115390 10834 115442 10846
rect 115390 10770 115442 10782
rect 116734 10834 116786 10846
rect 116734 10770 116786 10782
rect 37998 10722 38050 10734
rect 37998 10658 38050 10670
rect 47630 10722 47682 10734
rect 47630 10658 47682 10670
rect 51774 10722 51826 10734
rect 57486 10722 57538 10734
rect 53218 10670 53230 10722
rect 53282 10670 53294 10722
rect 51774 10658 51826 10670
rect 57486 10658 57538 10670
rect 73950 10722 74002 10734
rect 73950 10658 74002 10670
rect 74958 10722 75010 10734
rect 103518 10722 103570 10734
rect 83458 10670 83470 10722
rect 83522 10670 83534 10722
rect 74958 10658 75010 10670
rect 103518 10658 103570 10670
rect 104190 10722 104242 10734
rect 104190 10658 104242 10670
rect 105310 10722 105362 10734
rect 105310 10658 105362 10670
rect 57822 10610 57874 10622
rect 73390 10610 73442 10622
rect 37762 10558 37774 10610
rect 37826 10558 37838 10610
rect 42690 10558 42702 10610
rect 42754 10558 42766 10610
rect 47842 10558 47854 10610
rect 47906 10558 47918 10610
rect 52434 10558 52446 10610
rect 52498 10558 52510 10610
rect 61618 10558 61630 10610
rect 61682 10558 61694 10610
rect 62290 10558 62302 10610
rect 62354 10558 62366 10610
rect 68786 10558 68798 10610
rect 68850 10558 68862 10610
rect 72482 10558 72494 10610
rect 72546 10558 72558 10610
rect 57822 10546 57874 10558
rect 73390 10546 73442 10558
rect 74846 10610 74898 10622
rect 74846 10546 74898 10558
rect 75182 10610 75234 10622
rect 81790 10610 81842 10622
rect 79762 10558 79774 10610
rect 79826 10558 79838 10610
rect 82674 10558 82686 10610
rect 82738 10558 82750 10610
rect 86146 10558 86158 10610
rect 86210 10558 86222 10610
rect 88162 10558 88174 10610
rect 88226 10558 88238 10610
rect 92418 10558 92430 10610
rect 92482 10558 92494 10610
rect 100146 10558 100158 10610
rect 100210 10558 100222 10610
rect 109106 10558 109118 10610
rect 109170 10558 109182 10610
rect 75182 10546 75234 10558
rect 81790 10546 81842 10558
rect 38782 10498 38834 10510
rect 38782 10434 38834 10446
rect 39902 10498 39954 10510
rect 46062 10498 46114 10510
rect 43362 10446 43374 10498
rect 43426 10446 43438 10498
rect 45490 10446 45502 10498
rect 45554 10446 45566 10498
rect 39902 10434 39954 10446
rect 46062 10434 46114 10446
rect 47182 10498 47234 10510
rect 47182 10434 47234 10446
rect 49870 10498 49922 10510
rect 49870 10434 49922 10446
rect 50654 10498 50706 10510
rect 50654 10434 50706 10446
rect 51214 10498 51266 10510
rect 56478 10498 56530 10510
rect 55346 10446 55358 10498
rect 55410 10446 55422 10498
rect 51214 10434 51266 10446
rect 56478 10434 56530 10446
rect 58270 10498 58322 10510
rect 58270 10434 58322 10446
rect 58830 10498 58882 10510
rect 62862 10498 62914 10510
rect 59490 10446 59502 10498
rect 59554 10446 59566 10498
rect 58830 10434 58882 10446
rect 62862 10434 62914 10446
rect 63758 10498 63810 10510
rect 63758 10434 63810 10446
rect 64206 10498 64258 10510
rect 64206 10434 64258 10446
rect 64766 10498 64818 10510
rect 69694 10498 69746 10510
rect 76190 10498 76242 10510
rect 80446 10498 80498 10510
rect 65986 10446 65998 10498
rect 66050 10446 66062 10498
rect 68114 10446 68126 10498
rect 68178 10446 68190 10498
rect 71810 10446 71822 10498
rect 71874 10446 71886 10498
rect 79090 10446 79102 10498
rect 79154 10446 79166 10498
rect 64766 10434 64818 10446
rect 69694 10434 69746 10446
rect 76190 10434 76242 10446
rect 80446 10434 80498 10446
rect 81230 10498 81282 10510
rect 87054 10498 87106 10510
rect 85586 10446 85598 10498
rect 85650 10446 85662 10498
rect 81230 10434 81282 10446
rect 87054 10434 87106 10446
rect 87614 10498 87666 10510
rect 89518 10498 89570 10510
rect 96014 10498 96066 10510
rect 101950 10498 102002 10510
rect 88274 10446 88286 10498
rect 88338 10446 88350 10498
rect 91634 10446 91646 10498
rect 91698 10446 91710 10498
rect 97234 10446 97246 10498
rect 97298 10446 97310 10498
rect 99362 10446 99374 10498
rect 99426 10446 99438 10498
rect 87614 10434 87666 10446
rect 89518 10434 89570 10446
rect 96014 10434 96066 10446
rect 101950 10434 102002 10446
rect 102398 10498 102450 10510
rect 102398 10434 102450 10446
rect 102958 10498 103010 10510
rect 102958 10434 103010 10446
rect 106094 10498 106146 10510
rect 106094 10434 106146 10446
rect 106990 10498 107042 10510
rect 106990 10434 107042 10446
rect 107326 10498 107378 10510
rect 107326 10434 107378 10446
rect 108222 10498 108274 10510
rect 112030 10498 112082 10510
rect 109890 10446 109902 10498
rect 109954 10446 109966 10498
rect 108222 10434 108274 10446
rect 112030 10434 112082 10446
rect 113150 10498 113202 10510
rect 113150 10434 113202 10446
rect 113598 10498 113650 10510
rect 113598 10434 113650 10446
rect 113934 10498 113986 10510
rect 113934 10434 113986 10446
rect 114494 10498 114546 10510
rect 114494 10434 114546 10446
rect 115950 10498 116002 10510
rect 115950 10434 116002 10446
rect 117294 10498 117346 10510
rect 117294 10434 117346 10446
rect 117742 10498 117794 10510
rect 117742 10434 117794 10446
rect 118190 10498 118242 10510
rect 118190 10434 118242 10446
rect 51662 10386 51714 10398
rect 86494 10386 86546 10398
rect 58034 10334 58046 10386
rect 58098 10383 58110 10386
rect 58258 10383 58270 10386
rect 58098 10337 58270 10383
rect 58098 10334 58110 10337
rect 58258 10334 58270 10337
rect 58322 10383 58334 10386
rect 58706 10383 58718 10386
rect 58322 10337 58718 10383
rect 58322 10334 58334 10337
rect 58706 10334 58718 10337
rect 58770 10334 58782 10386
rect 51662 10322 51714 10334
rect 86494 10322 86546 10334
rect 88510 10386 88562 10398
rect 104414 10386 104466 10398
rect 101266 10334 101278 10386
rect 101330 10383 101342 10386
rect 101938 10383 101950 10386
rect 101330 10337 101950 10383
rect 101330 10334 101342 10337
rect 101938 10334 101950 10337
rect 102002 10334 102014 10386
rect 88510 10322 88562 10334
rect 104414 10322 104466 10334
rect 105534 10386 105586 10398
rect 106530 10334 106542 10386
rect 106594 10383 106606 10386
rect 107314 10383 107326 10386
rect 106594 10337 107326 10383
rect 106594 10334 106606 10337
rect 107314 10334 107326 10337
rect 107378 10334 107390 10386
rect 105534 10322 105586 10334
rect 1344 10218 178640 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 96638 10218
rect 96690 10166 96742 10218
rect 96794 10166 96846 10218
rect 96898 10166 127358 10218
rect 127410 10166 127462 10218
rect 127514 10166 127566 10218
rect 127618 10166 158078 10218
rect 158130 10166 158182 10218
rect 158234 10166 158286 10218
rect 158338 10166 178640 10218
rect 1344 10132 178640 10166
rect 51774 10050 51826 10062
rect 51774 9986 51826 9998
rect 52670 10050 52722 10062
rect 52670 9986 52722 9998
rect 54350 10050 54402 10062
rect 54350 9986 54402 9998
rect 54686 10050 54738 10062
rect 83582 10050 83634 10062
rect 95454 10050 95506 10062
rect 118190 10050 118242 10062
rect 61730 9998 61742 10050
rect 61794 10047 61806 10050
rect 62066 10047 62078 10050
rect 61794 10001 62078 10047
rect 61794 9998 61806 10001
rect 62066 9998 62078 10001
rect 62130 9998 62142 10050
rect 86930 9998 86942 10050
rect 86994 10047 87006 10050
rect 87154 10047 87166 10050
rect 86994 10001 87166 10047
rect 86994 9998 87006 10001
rect 87154 9998 87166 10001
rect 87218 9998 87230 10050
rect 104402 9998 104414 10050
rect 104466 10047 104478 10050
rect 104626 10047 104638 10050
rect 104466 10001 104638 10047
rect 104466 9998 104478 10001
rect 104626 9998 104638 10001
rect 104690 9998 104702 10050
rect 106530 9998 106542 10050
rect 106594 10047 106606 10050
rect 106978 10047 106990 10050
rect 106594 10001 106990 10047
rect 106594 9998 106606 10001
rect 106978 9998 106990 10001
rect 107042 9998 107054 10050
rect 114818 9998 114830 10050
rect 114882 10047 114894 10050
rect 115490 10047 115502 10050
rect 114882 10001 115502 10047
rect 114882 9998 114894 10001
rect 115490 9998 115502 10001
rect 115554 9998 115566 10050
rect 54686 9986 54738 9998
rect 83582 9986 83634 9998
rect 95454 9986 95506 9998
rect 118190 9986 118242 9998
rect 119086 10050 119138 10062
rect 119086 9986 119138 9998
rect 40910 9938 40962 9950
rect 33506 9886 33518 9938
rect 33570 9886 33582 9938
rect 38322 9886 38334 9938
rect 38386 9886 38398 9938
rect 40450 9886 40462 9938
rect 40514 9886 40526 9938
rect 40910 9874 40962 9886
rect 43150 9938 43202 9950
rect 50878 9938 50930 9950
rect 47394 9886 47406 9938
rect 47458 9886 47470 9938
rect 49522 9886 49534 9938
rect 49586 9886 49598 9938
rect 43150 9874 43202 9886
rect 50878 9874 50930 9886
rect 53678 9938 53730 9950
rect 61742 9938 61794 9950
rect 56914 9886 56926 9938
rect 56978 9886 56990 9938
rect 59042 9886 59054 9938
rect 59106 9886 59118 9938
rect 53678 9874 53730 9886
rect 61742 9874 61794 9886
rect 62190 9938 62242 9950
rect 62190 9874 62242 9886
rect 63422 9938 63474 9950
rect 63422 9874 63474 9886
rect 63982 9938 64034 9950
rect 63982 9874 64034 9886
rect 64766 9938 64818 9950
rect 75294 9938 75346 9950
rect 78654 9938 78706 9950
rect 73826 9886 73838 9938
rect 73890 9886 73902 9938
rect 76178 9886 76190 9938
rect 76242 9886 76254 9938
rect 64766 9874 64818 9886
rect 75294 9874 75346 9886
rect 78654 9874 78706 9886
rect 84590 9938 84642 9950
rect 84590 9874 84642 9886
rect 85822 9938 85874 9950
rect 85822 9874 85874 9886
rect 86942 9938 86994 9950
rect 86942 9874 86994 9886
rect 100270 9938 100322 9950
rect 100270 9874 100322 9886
rect 103294 9938 103346 9950
rect 103294 9874 103346 9886
rect 103630 9938 103682 9950
rect 103630 9874 103682 9886
rect 104078 9938 104130 9950
rect 104078 9874 104130 9886
rect 105198 9938 105250 9950
rect 105198 9874 105250 9886
rect 106430 9938 106482 9950
rect 106430 9874 106482 9886
rect 106990 9938 107042 9950
rect 106990 9874 107042 9886
rect 108334 9938 108386 9950
rect 108334 9874 108386 9886
rect 112142 9938 112194 9950
rect 112142 9874 112194 9886
rect 113262 9938 113314 9950
rect 113262 9874 113314 9886
rect 114158 9938 114210 9950
rect 114158 9874 114210 9886
rect 116062 9938 116114 9950
rect 116062 9874 116114 9886
rect 60174 9826 60226 9838
rect 81006 9826 81058 9838
rect 30706 9774 30718 9826
rect 30770 9774 30782 9826
rect 37650 9774 37662 9826
rect 37714 9774 37726 9826
rect 45602 9774 45614 9826
rect 45666 9774 45678 9826
rect 46722 9774 46734 9826
rect 46786 9774 46798 9826
rect 51426 9774 51438 9826
rect 51490 9774 51502 9826
rect 52322 9774 52334 9826
rect 52386 9774 52398 9826
rect 55458 9774 55470 9826
rect 55522 9774 55534 9826
rect 56130 9774 56142 9826
rect 56194 9774 56206 9826
rect 68338 9774 68350 9826
rect 68402 9774 68414 9826
rect 69346 9774 69358 9826
rect 69410 9774 69422 9826
rect 77746 9774 77758 9826
rect 77810 9774 77822 9826
rect 60174 9762 60226 9774
rect 81006 9762 81058 9774
rect 81454 9826 81506 9838
rect 81454 9762 81506 9774
rect 82238 9826 82290 9838
rect 98142 9826 98194 9838
rect 88274 9774 88286 9826
rect 88338 9774 88350 9826
rect 82238 9762 82290 9774
rect 98142 9762 98194 9774
rect 98814 9826 98866 9838
rect 102734 9826 102786 9838
rect 117182 9826 117234 9838
rect 99138 9774 99150 9826
rect 99202 9774 99214 9826
rect 109218 9774 109230 9826
rect 109282 9774 109294 9826
rect 98814 9762 98866 9774
rect 102734 9762 102786 9774
rect 117182 9762 117234 9774
rect 36542 9714 36594 9726
rect 31378 9662 31390 9714
rect 31442 9662 31454 9714
rect 36542 9650 36594 9662
rect 43710 9714 43762 9726
rect 43710 9650 43762 9662
rect 44046 9714 44098 9726
rect 44046 9650 44098 9662
rect 50430 9714 50482 9726
rect 60510 9714 60562 9726
rect 75182 9714 75234 9726
rect 55234 9662 55246 9714
rect 55298 9662 55310 9714
rect 67666 9662 67678 9714
rect 67730 9662 67742 9714
rect 50430 9650 50482 9662
rect 60510 9650 60562 9662
rect 75182 9650 75234 9662
rect 76526 9714 76578 9726
rect 76526 9650 76578 9662
rect 78766 9714 78818 9726
rect 78766 9650 78818 9662
rect 79214 9714 79266 9726
rect 79214 9650 79266 9662
rect 83918 9714 83970 9726
rect 83918 9650 83970 9662
rect 87614 9714 87666 9726
rect 87614 9650 87666 9662
rect 87726 9714 87778 9726
rect 95790 9714 95842 9726
rect 89058 9662 89070 9714
rect 89122 9662 89134 9714
rect 87726 9650 87778 9662
rect 95790 9650 95842 9662
rect 96574 9714 96626 9726
rect 96574 9650 96626 9662
rect 96910 9714 96962 9726
rect 96910 9650 96962 9662
rect 97694 9714 97746 9726
rect 97694 9650 97746 9662
rect 98366 9714 98418 9726
rect 98366 9650 98418 9662
rect 101054 9714 101106 9726
rect 101054 9650 101106 9662
rect 102398 9714 102450 9726
rect 117070 9714 117122 9726
rect 110002 9662 110014 9714
rect 110066 9662 110078 9714
rect 102398 9650 102450 9662
rect 117070 9650 117122 9662
rect 117294 9714 117346 9726
rect 117294 9650 117346 9662
rect 118526 9714 118578 9726
rect 118526 9650 118578 9662
rect 119198 9714 119250 9726
rect 119198 9650 119250 9662
rect 119422 9714 119474 9726
rect 119422 9650 119474 9662
rect 33966 9602 34018 9614
rect 33966 9538 34018 9550
rect 35198 9602 35250 9614
rect 35198 9538 35250 9550
rect 36206 9602 36258 9614
rect 36206 9538 36258 9550
rect 41470 9602 41522 9614
rect 41470 9538 41522 9550
rect 42142 9602 42194 9614
rect 42142 9538 42194 9550
rect 42590 9602 42642 9614
rect 42590 9538 42642 9550
rect 44830 9602 44882 9614
rect 44830 9538 44882 9550
rect 45838 9602 45890 9614
rect 45838 9538 45890 9550
rect 50094 9602 50146 9614
rect 50094 9538 50146 9550
rect 51662 9602 51714 9614
rect 51662 9538 51714 9550
rect 52558 9602 52610 9614
rect 52558 9538 52610 9550
rect 59614 9602 59666 9614
rect 59614 9538 59666 9550
rect 62526 9602 62578 9614
rect 62526 9538 62578 9550
rect 62974 9602 63026 9614
rect 62974 9538 63026 9550
rect 64318 9602 64370 9614
rect 75406 9602 75458 9614
rect 65426 9550 65438 9602
rect 65490 9550 65502 9602
rect 64318 9538 64370 9550
rect 75406 9538 75458 9550
rect 76302 9602 76354 9614
rect 76302 9538 76354 9550
rect 77534 9602 77586 9614
rect 77534 9538 77586 9550
rect 78542 9602 78594 9614
rect 78542 9538 78594 9550
rect 79662 9602 79714 9614
rect 79662 9538 79714 9550
rect 80110 9602 80162 9614
rect 80110 9538 80162 9550
rect 80670 9602 80722 9614
rect 80670 9538 80722 9550
rect 82574 9602 82626 9614
rect 82574 9538 82626 9550
rect 83134 9602 83186 9614
rect 83134 9538 83186 9550
rect 83694 9602 83746 9614
rect 83694 9538 83746 9550
rect 85486 9602 85538 9614
rect 85486 9538 85538 9550
rect 86494 9602 86546 9614
rect 86494 9538 86546 9550
rect 87502 9602 87554 9614
rect 95006 9602 95058 9614
rect 91298 9550 91310 9602
rect 91362 9550 91374 9602
rect 87502 9538 87554 9550
rect 95006 9538 95058 9550
rect 95566 9602 95618 9614
rect 95566 9538 95618 9550
rect 97582 9602 97634 9614
rect 97582 9538 97634 9550
rect 97918 9602 97970 9614
rect 97918 9538 97970 9550
rect 99374 9602 99426 9614
rect 99374 9538 99426 9550
rect 99486 9602 99538 9614
rect 99486 9538 99538 9550
rect 99822 9602 99874 9614
rect 99822 9538 99874 9550
rect 101502 9602 101554 9614
rect 101502 9538 101554 9550
rect 104638 9602 104690 9614
rect 104638 9538 104690 9550
rect 105534 9602 105586 9614
rect 105534 9538 105586 9550
rect 105982 9602 106034 9614
rect 105982 9538 106034 9550
rect 107438 9602 107490 9614
rect 107438 9538 107490 9550
rect 107886 9602 107938 9614
rect 107886 9538 107938 9550
rect 112814 9602 112866 9614
rect 112814 9538 112866 9550
rect 113710 9602 113762 9614
rect 113710 9538 113762 9550
rect 114718 9602 114770 9614
rect 114718 9538 114770 9550
rect 115054 9602 115106 9614
rect 115054 9538 115106 9550
rect 115502 9602 115554 9614
rect 115502 9538 115554 9550
rect 118302 9602 118354 9614
rect 118302 9538 118354 9550
rect 119870 9602 119922 9614
rect 119870 9538 119922 9550
rect 1344 9434 178640 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 81278 9434
rect 81330 9382 81382 9434
rect 81434 9382 81486 9434
rect 81538 9382 111998 9434
rect 112050 9382 112102 9434
rect 112154 9382 112206 9434
rect 112258 9382 142718 9434
rect 142770 9382 142822 9434
rect 142874 9382 142926 9434
rect 142978 9382 173438 9434
rect 173490 9382 173542 9434
rect 173594 9382 173646 9434
rect 173698 9382 178640 9434
rect 1344 9348 178640 9382
rect 31838 9266 31890 9278
rect 31838 9202 31890 9214
rect 32846 9266 32898 9278
rect 32846 9202 32898 9214
rect 35422 9266 35474 9278
rect 35422 9202 35474 9214
rect 36990 9266 37042 9278
rect 36990 9202 37042 9214
rect 41470 9266 41522 9278
rect 41470 9202 41522 9214
rect 41918 9266 41970 9278
rect 41918 9202 41970 9214
rect 42590 9266 42642 9278
rect 42590 9202 42642 9214
rect 43038 9266 43090 9278
rect 43038 9202 43090 9214
rect 43486 9266 43538 9278
rect 43486 9202 43538 9214
rect 44606 9266 44658 9278
rect 44606 9202 44658 9214
rect 46846 9266 46898 9278
rect 46846 9202 46898 9214
rect 47518 9266 47570 9278
rect 47518 9202 47570 9214
rect 55694 9266 55746 9278
rect 55694 9202 55746 9214
rect 57934 9266 57986 9278
rect 57934 9202 57986 9214
rect 65438 9266 65490 9278
rect 65438 9202 65490 9214
rect 65774 9266 65826 9278
rect 65774 9202 65826 9214
rect 66222 9266 66274 9278
rect 66222 9202 66274 9214
rect 66894 9266 66946 9278
rect 66894 9202 66946 9214
rect 67790 9266 67842 9278
rect 67790 9202 67842 9214
rect 67902 9266 67954 9278
rect 67902 9202 67954 9214
rect 68686 9266 68738 9278
rect 68686 9202 68738 9214
rect 73726 9266 73778 9278
rect 73726 9202 73778 9214
rect 74622 9266 74674 9278
rect 74622 9202 74674 9214
rect 79662 9266 79714 9278
rect 79662 9202 79714 9214
rect 80558 9266 80610 9278
rect 80558 9202 80610 9214
rect 81566 9266 81618 9278
rect 81566 9202 81618 9214
rect 88062 9266 88114 9278
rect 94670 9266 94722 9278
rect 90178 9214 90190 9266
rect 90242 9214 90254 9266
rect 88062 9202 88114 9214
rect 94670 9202 94722 9214
rect 96238 9266 96290 9278
rect 96238 9202 96290 9214
rect 99822 9266 99874 9278
rect 99822 9202 99874 9214
rect 100494 9266 100546 9278
rect 100494 9202 100546 9214
rect 100942 9266 100994 9278
rect 100942 9202 100994 9214
rect 108558 9266 108610 9278
rect 114382 9266 114434 9278
rect 113698 9214 113710 9266
rect 113762 9263 113774 9266
rect 113762 9217 113871 9263
rect 113762 9214 113774 9217
rect 108558 9202 108610 9214
rect 46510 9154 46562 9166
rect 55358 9154 55410 9166
rect 59614 9154 59666 9166
rect 89406 9154 89458 9166
rect 95118 9154 95170 9166
rect 34626 9102 34638 9154
rect 34690 9102 34702 9154
rect 45490 9102 45502 9154
rect 45554 9102 45566 9154
rect 48626 9102 48638 9154
rect 48690 9102 48702 9154
rect 53554 9102 53566 9154
rect 53618 9102 53630 9154
rect 58594 9102 58606 9154
rect 58658 9102 58670 9154
rect 58818 9102 58830 9154
rect 58882 9102 58894 9154
rect 71810 9102 71822 9154
rect 71874 9102 71886 9154
rect 76066 9102 76078 9154
rect 76130 9102 76142 9154
rect 94770 9102 94782 9154
rect 94834 9151 94846 9154
rect 94994 9151 95006 9154
rect 94834 9105 95006 9151
rect 94834 9102 94846 9105
rect 94994 9102 95006 9105
rect 95058 9102 95070 9154
rect 46510 9090 46562 9102
rect 55358 9090 55410 9102
rect 59614 9090 59666 9102
rect 89406 9090 89458 9102
rect 95118 9090 95170 9102
rect 96462 9154 96514 9166
rect 96462 9090 96514 9102
rect 97358 9154 97410 9166
rect 97358 9090 97410 9102
rect 99486 9154 99538 9166
rect 99486 9090 99538 9102
rect 113038 9154 113090 9166
rect 113038 9090 113090 9102
rect 32174 9042 32226 9054
rect 32174 8978 32226 8990
rect 33742 9042 33794 9054
rect 33742 8978 33794 8990
rect 34078 9042 34130 9054
rect 44942 9042 44994 9054
rect 47854 9042 47906 9054
rect 56142 9042 56194 9054
rect 34514 8990 34526 9042
rect 34578 8990 34590 9042
rect 37986 8990 37998 9042
rect 38050 8990 38062 9042
rect 45714 8990 45726 9042
rect 45778 8990 45790 9042
rect 48402 8990 48414 9042
rect 48466 8990 48478 9042
rect 50306 8990 50318 9042
rect 50370 8990 50382 9042
rect 34078 8978 34130 8990
rect 44942 8978 44994 8990
rect 47854 8978 47906 8990
rect 56142 8978 56194 8990
rect 56702 9042 56754 9054
rect 74510 9042 74562 9054
rect 83022 9042 83074 9054
rect 89294 9042 89346 9054
rect 60610 8990 60622 9042
rect 60674 8990 60686 9042
rect 64418 8990 64430 9042
rect 64482 8990 64494 9042
rect 72482 8990 72494 9042
rect 72546 8990 72558 9042
rect 75394 8990 75406 9042
rect 75458 8990 75470 9042
rect 82114 8990 82126 9042
rect 82178 8990 82190 9042
rect 86482 8990 86494 9042
rect 86546 8990 86558 9042
rect 56702 8978 56754 8990
rect 74510 8978 74562 8990
rect 83022 8978 83074 8990
rect 89294 8978 89346 8990
rect 89630 9042 89682 9054
rect 95902 9042 95954 9054
rect 98814 9042 98866 9054
rect 93202 8990 93214 9042
rect 93266 8990 93278 9042
rect 98354 8990 98366 9042
rect 98418 8990 98430 9042
rect 89630 8978 89682 8990
rect 95902 8978 95954 8990
rect 98814 8978 98866 8990
rect 99710 9042 99762 9054
rect 99710 8978 99762 8990
rect 100158 9042 100210 9054
rect 104290 8990 104302 9042
rect 104354 8990 104366 9042
rect 105186 8990 105198 9042
rect 105250 8990 105262 9042
rect 109106 8990 109118 9042
rect 109170 8990 109182 9042
rect 100158 8978 100210 8990
rect 35870 8930 35922 8942
rect 35870 8866 35922 8878
rect 36318 8930 36370 8942
rect 36318 8866 36370 8878
rect 37438 8930 37490 8942
rect 44046 8930 44098 8942
rect 38658 8878 38670 8930
rect 38722 8878 38734 8930
rect 40786 8878 40798 8930
rect 40850 8878 40862 8930
rect 37438 8866 37490 8878
rect 44046 8866 44098 8878
rect 58270 8930 58322 8942
rect 64206 8930 64258 8942
rect 69694 8930 69746 8942
rect 78766 8930 78818 8942
rect 61282 8878 61294 8930
rect 61346 8878 61358 8930
rect 63410 8878 63422 8930
rect 63474 8878 63486 8930
rect 66770 8878 66782 8930
rect 66834 8878 66846 8930
rect 68562 8878 68574 8930
rect 68626 8878 68638 8930
rect 73602 8878 73614 8930
rect 73666 8878 73678 8930
rect 78194 8878 78206 8930
rect 78258 8878 78270 8930
rect 58270 8866 58322 8878
rect 64206 8866 64258 8878
rect 69694 8866 69746 8878
rect 78766 8866 78818 8878
rect 80110 8930 80162 8942
rect 86942 8930 86994 8942
rect 83570 8878 83582 8930
rect 83634 8878 83646 8930
rect 85698 8878 85710 8930
rect 85762 8878 85774 8930
rect 80110 8866 80162 8878
rect 86942 8866 86994 8878
rect 87614 8930 87666 8942
rect 87614 8866 87666 8878
rect 88510 8930 88562 8942
rect 94222 8930 94274 8942
rect 92418 8878 92430 8930
rect 92482 8878 92494 8930
rect 88510 8866 88562 8878
rect 94222 8866 94274 8878
rect 98926 8930 98978 8942
rect 113486 8930 113538 8942
rect 101490 8878 101502 8930
rect 101554 8878 101566 8930
rect 103618 8878 103630 8930
rect 103682 8878 103694 8930
rect 105970 8878 105982 8930
rect 106034 8878 106046 8930
rect 108098 8878 108110 8930
rect 108162 8878 108174 8930
rect 109890 8878 109902 8930
rect 109954 8878 109966 8930
rect 112018 8878 112030 8930
rect 112082 8878 112094 8930
rect 98926 8866 98978 8878
rect 113486 8866 113538 8878
rect 64094 8818 64146 8830
rect 35746 8766 35758 8818
rect 35810 8815 35822 8818
rect 36306 8815 36318 8818
rect 35810 8769 36318 8815
rect 35810 8766 35822 8769
rect 36306 8766 36318 8769
rect 36370 8766 36382 8818
rect 64094 8754 64146 8766
rect 67118 8818 67170 8830
rect 67118 8754 67170 8766
rect 68014 8818 68066 8830
rect 68014 8754 68066 8766
rect 68910 8818 68962 8830
rect 68910 8754 68962 8766
rect 73950 8818 74002 8830
rect 73950 8754 74002 8766
rect 74622 8818 74674 8830
rect 74622 8754 74674 8766
rect 78878 8818 78930 8830
rect 78878 8754 78930 8766
rect 82126 8818 82178 8830
rect 82126 8754 82178 8766
rect 82462 8818 82514 8830
rect 82462 8754 82514 8766
rect 95230 8818 95282 8830
rect 95230 8754 95282 8766
rect 96574 8818 96626 8830
rect 96574 8754 96626 8766
rect 97246 8818 97298 8830
rect 113825 8818 113871 9217
rect 114382 9202 114434 9214
rect 114830 9266 114882 9278
rect 114830 9202 114882 9214
rect 116622 9266 116674 9278
rect 116622 9202 116674 9214
rect 118638 9266 118690 9278
rect 118638 9202 118690 9214
rect 120990 9266 121042 9278
rect 120990 9202 121042 9214
rect 121886 9266 121938 9278
rect 121886 9202 121938 9214
rect 115390 9154 115442 9166
rect 115390 9090 115442 9102
rect 115726 9154 115778 9166
rect 115726 9090 115778 9102
rect 116286 9154 116338 9166
rect 116286 9090 116338 9102
rect 117182 9154 117234 9166
rect 117182 9090 117234 9102
rect 117518 9154 117570 9166
rect 117518 9090 117570 9102
rect 114046 9042 114098 9054
rect 121550 9042 121602 9054
rect 118402 8990 118414 9042
rect 118466 8990 118478 9042
rect 114046 8978 114098 8990
rect 121550 8978 121602 8990
rect 119198 8930 119250 8942
rect 119198 8866 119250 8878
rect 119646 8930 119698 8942
rect 119646 8866 119698 8878
rect 120094 8930 120146 8942
rect 120094 8866 120146 8878
rect 118750 8818 118802 8830
rect 113810 8766 113822 8818
rect 113874 8766 113886 8818
rect 119522 8766 119534 8818
rect 119586 8815 119598 8818
rect 120082 8815 120094 8818
rect 119586 8769 120094 8815
rect 119586 8766 119598 8769
rect 120082 8766 120094 8769
rect 120146 8766 120158 8818
rect 97246 8754 97298 8766
rect 118750 8754 118802 8766
rect 1344 8650 178640 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 96638 8650
rect 96690 8598 96742 8650
rect 96794 8598 96846 8650
rect 96898 8598 127358 8650
rect 127410 8598 127462 8650
rect 127514 8598 127566 8650
rect 127618 8598 158078 8650
rect 158130 8598 158182 8650
rect 158234 8598 158286 8650
rect 158338 8598 178640 8650
rect 1344 8564 178640 8598
rect 38222 8482 38274 8494
rect 94782 8482 94834 8494
rect 42466 8430 42478 8482
rect 42530 8479 42542 8482
rect 43138 8479 43150 8482
rect 42530 8433 43150 8479
rect 42530 8430 42542 8433
rect 43138 8430 43150 8433
rect 43202 8430 43214 8482
rect 59714 8430 59726 8482
rect 59778 8479 59790 8482
rect 60050 8479 60062 8482
rect 59778 8433 60062 8479
rect 59778 8430 59790 8433
rect 60050 8430 60062 8433
rect 60114 8430 60126 8482
rect 38222 8418 38274 8430
rect 94782 8418 94834 8430
rect 98814 8482 98866 8494
rect 100370 8479 100382 8482
rect 98814 8418 98866 8430
rect 100049 8433 100382 8479
rect 37886 8370 37938 8382
rect 33618 8318 33630 8370
rect 33682 8318 33694 8370
rect 37886 8306 37938 8318
rect 40126 8370 40178 8382
rect 40126 8306 40178 8318
rect 43038 8370 43090 8382
rect 43038 8306 43090 8318
rect 43934 8370 43986 8382
rect 60174 8370 60226 8382
rect 48178 8318 48190 8370
rect 48242 8318 48254 8370
rect 50306 8318 50318 8370
rect 50370 8318 50382 8370
rect 55234 8318 55246 8370
rect 55298 8318 55310 8370
rect 43934 8306 43986 8318
rect 60174 8306 60226 8318
rect 68238 8370 68290 8382
rect 83694 8370 83746 8382
rect 68562 8318 68574 8370
rect 68626 8318 68638 8370
rect 73490 8318 73502 8370
rect 73554 8318 73566 8370
rect 78530 8318 78542 8370
rect 78594 8318 78606 8370
rect 82450 8318 82462 8370
rect 82514 8318 82526 8370
rect 68238 8306 68290 8318
rect 83694 8306 83746 8318
rect 85710 8370 85762 8382
rect 85710 8306 85762 8318
rect 86270 8370 86322 8382
rect 91870 8370 91922 8382
rect 90290 8318 90302 8370
rect 90354 8318 90366 8370
rect 86270 8306 86322 8318
rect 91870 8306 91922 8318
rect 92430 8370 92482 8382
rect 92430 8306 92482 8318
rect 93774 8370 93826 8382
rect 93774 8306 93826 8318
rect 94222 8370 94274 8382
rect 94222 8306 94274 8318
rect 95342 8370 95394 8382
rect 100049 8370 100095 8433
rect 100370 8430 100382 8433
rect 100434 8430 100446 8482
rect 100158 8370 100210 8382
rect 100034 8318 100046 8370
rect 100098 8318 100110 8370
rect 95342 8306 95394 8318
rect 100158 8306 100210 8318
rect 101838 8370 101890 8382
rect 101838 8306 101890 8318
rect 105198 8370 105250 8382
rect 105198 8306 105250 8318
rect 113262 8370 113314 8382
rect 113262 8306 113314 8318
rect 117518 8370 117570 8382
rect 117518 8306 117570 8318
rect 123454 8370 123506 8382
rect 123454 8306 123506 8318
rect 138798 8370 138850 8382
rect 138798 8306 138850 8318
rect 35086 8258 35138 8270
rect 45502 8258 45554 8270
rect 51886 8258 51938 8270
rect 30706 8206 30718 8258
rect 30770 8206 30782 8258
rect 38882 8206 38894 8258
rect 38946 8206 38958 8258
rect 50978 8206 50990 8258
rect 51042 8206 51054 8258
rect 35086 8194 35138 8206
rect 45502 8194 45554 8206
rect 51886 8194 51938 8206
rect 52110 8258 52162 8270
rect 52110 8194 52162 8206
rect 52446 8258 52498 8270
rect 52446 8194 52498 8206
rect 53342 8258 53394 8270
rect 53342 8194 53394 8206
rect 54014 8258 54066 8270
rect 54014 8194 54066 8206
rect 54798 8258 54850 8270
rect 54798 8194 54850 8206
rect 59278 8258 59330 8270
rect 67342 8258 67394 8270
rect 75406 8258 75458 8270
rect 78990 8258 79042 8270
rect 61394 8206 61406 8258
rect 61458 8206 61470 8258
rect 69346 8206 69358 8258
rect 69410 8206 69422 8258
rect 77410 8206 77422 8258
rect 77474 8206 77486 8258
rect 59278 8194 59330 8206
rect 67342 8194 67394 8206
rect 75406 8194 75458 8206
rect 78990 8194 79042 8206
rect 80670 8258 80722 8270
rect 80670 8194 80722 8206
rect 80894 8258 80946 8270
rect 80894 8194 80946 8206
rect 81118 8258 81170 8270
rect 84254 8258 84306 8270
rect 82562 8206 82574 8258
rect 82626 8206 82638 8258
rect 81118 8194 81170 8206
rect 84254 8194 84306 8206
rect 84590 8258 84642 8270
rect 84590 8194 84642 8206
rect 85486 8258 85538 8270
rect 85486 8194 85538 8206
rect 87278 8258 87330 8270
rect 87278 8194 87330 8206
rect 87502 8258 87554 8270
rect 94894 8258 94946 8270
rect 90178 8206 90190 8258
rect 90242 8206 90254 8258
rect 91634 8206 91646 8258
rect 91698 8206 91710 8258
rect 87502 8194 87554 8206
rect 94894 8194 94946 8206
rect 95566 8258 95618 8270
rect 95566 8194 95618 8206
rect 96350 8258 96402 8270
rect 96350 8194 96402 8206
rect 97806 8258 97858 8270
rect 97806 8194 97858 8206
rect 98590 8258 98642 8270
rect 98590 8194 98642 8206
rect 99150 8258 99202 8270
rect 101390 8258 101442 8270
rect 99474 8206 99486 8258
rect 99538 8206 99550 8258
rect 99150 8194 99202 8206
rect 101390 8194 101442 8206
rect 102846 8258 102898 8270
rect 104414 8258 104466 8270
rect 103730 8206 103742 8258
rect 103794 8206 103806 8258
rect 102846 8194 102898 8206
rect 104414 8194 104466 8206
rect 108334 8258 108386 8270
rect 116062 8258 116114 8270
rect 109330 8206 109342 8258
rect 109394 8206 109406 8258
rect 114930 8206 114942 8258
rect 114994 8206 115006 8258
rect 108334 8194 108386 8206
rect 116062 8194 116114 8206
rect 116958 8258 117010 8270
rect 116958 8194 117010 8206
rect 119646 8258 119698 8270
rect 119646 8194 119698 8206
rect 119758 8258 119810 8270
rect 119758 8194 119810 8206
rect 120654 8258 120706 8270
rect 120654 8194 120706 8206
rect 19630 8146 19682 8158
rect 19630 8082 19682 8094
rect 27134 8146 27186 8158
rect 36430 8146 36482 8158
rect 46398 8146 46450 8158
rect 31490 8094 31502 8146
rect 31554 8094 31566 8146
rect 34290 8094 34302 8146
rect 34354 8094 34366 8146
rect 34738 8094 34750 8146
rect 34802 8094 34814 8146
rect 38994 8094 39006 8146
rect 39058 8094 39070 8146
rect 40338 8094 40350 8146
rect 40402 8094 40414 8146
rect 40786 8094 40798 8146
rect 40850 8094 40862 8146
rect 27134 8082 27186 8094
rect 36430 8082 36482 8094
rect 46398 8082 46450 8094
rect 46734 8146 46786 8158
rect 46734 8082 46786 8094
rect 47294 8146 47346 8158
rect 47294 8082 47346 8094
rect 53790 8146 53842 8158
rect 53790 8082 53842 8094
rect 56254 8146 56306 8158
rect 56254 8082 56306 8094
rect 57486 8146 57538 8158
rect 57486 8082 57538 8094
rect 57822 8146 57874 8158
rect 75518 8146 75570 8158
rect 76526 8146 76578 8158
rect 66434 8094 66446 8146
rect 66498 8094 66510 8146
rect 76178 8094 76190 8146
rect 76242 8094 76254 8146
rect 57822 8082 57874 8094
rect 75518 8082 75570 8094
rect 76526 8082 76578 8094
rect 78206 8146 78258 8158
rect 78206 8082 78258 8094
rect 78430 8146 78482 8158
rect 78430 8082 78482 8094
rect 79326 8146 79378 8158
rect 79326 8082 79378 8094
rect 79886 8146 79938 8158
rect 79886 8082 79938 8094
rect 81342 8146 81394 8158
rect 81342 8082 81394 8094
rect 83246 8146 83298 8158
rect 83246 8082 83298 8094
rect 85262 8146 85314 8158
rect 85262 8082 85314 8094
rect 85822 8146 85874 8158
rect 85822 8082 85874 8094
rect 86718 8146 86770 8158
rect 88734 8146 88786 8158
rect 87826 8094 87838 8146
rect 87890 8094 87902 8146
rect 86718 8082 86770 8094
rect 88734 8082 88786 8094
rect 91086 8146 91138 8158
rect 91086 8082 91138 8094
rect 91982 8146 92034 8158
rect 91982 8082 92034 8094
rect 96686 8146 96738 8158
rect 96686 8082 96738 8094
rect 98030 8146 98082 8158
rect 98030 8082 98082 8094
rect 98142 8146 98194 8158
rect 98142 8082 98194 8094
rect 99710 8146 99762 8158
rect 99710 8082 99762 8094
rect 99822 8146 99874 8158
rect 99822 8082 99874 8094
rect 101614 8146 101666 8158
rect 101614 8082 101666 8094
rect 101950 8146 102002 8158
rect 101950 8082 102002 8094
rect 103966 8146 104018 8158
rect 103966 8082 104018 8094
rect 105310 8146 105362 8158
rect 105310 8082 105362 8094
rect 107214 8146 107266 8158
rect 113710 8146 113762 8158
rect 110002 8094 110014 8146
rect 110066 8094 110078 8146
rect 107214 8082 107266 8094
rect 113710 8082 113762 8094
rect 119534 8146 119586 8158
rect 119534 8082 119586 8094
rect 19294 8034 19346 8046
rect 19294 7970 19346 7982
rect 26798 8034 26850 8046
rect 26798 7970 26850 7982
rect 27806 8034 27858 8046
rect 27806 7970 27858 7982
rect 28814 8034 28866 8046
rect 28814 7970 28866 7982
rect 29598 8034 29650 8046
rect 29598 7970 29650 7982
rect 35422 8034 35474 8046
rect 35422 7970 35474 7982
rect 36878 8034 36930 8046
rect 36878 7970 36930 7982
rect 39790 8034 39842 8046
rect 39790 7970 39842 7982
rect 41806 8034 41858 8046
rect 41806 7970 41858 7982
rect 42254 8034 42306 8046
rect 42254 7970 42306 7982
rect 42590 8034 42642 8046
rect 42590 7970 42642 7982
rect 43710 8034 43762 8046
rect 43710 7970 43762 7982
rect 43822 8034 43874 8046
rect 43822 7970 43874 7982
rect 44830 8034 44882 8046
rect 44830 7970 44882 7982
rect 45838 8034 45890 8046
rect 45838 7970 45890 7982
rect 47630 8034 47682 8046
rect 47630 7970 47682 7982
rect 52334 8034 52386 8046
rect 52334 7970 52386 7982
rect 53566 8034 53618 8046
rect 53566 7970 53618 7982
rect 55918 8034 55970 8046
rect 55918 7970 55970 7982
rect 57038 8034 57090 8046
rect 57038 7970 57090 7982
rect 58382 8034 58434 8046
rect 58382 7970 58434 7982
rect 58942 8034 58994 8046
rect 58942 7970 58994 7982
rect 59726 8034 59778 8046
rect 59726 7970 59778 7982
rect 60734 8034 60786 8046
rect 60734 7970 60786 7982
rect 67678 8034 67730 8046
rect 67678 7970 67730 7982
rect 75742 8034 75794 8046
rect 75742 7970 75794 7982
rect 77646 8034 77698 8046
rect 77646 7970 77698 7982
rect 79214 8034 79266 8046
rect 79214 7970 79266 7982
rect 80222 8034 80274 8046
rect 80222 7970 80274 7982
rect 84366 8034 84418 8046
rect 84366 7970 84418 7982
rect 88398 8034 88450 8046
rect 88398 7970 88450 7982
rect 89406 8034 89458 8046
rect 89406 7970 89458 7982
rect 93102 8034 93154 8046
rect 93102 7970 93154 7982
rect 95678 8034 95730 8046
rect 95678 7970 95730 7982
rect 96238 8034 96290 8046
rect 96238 7970 96290 7982
rect 96462 8034 96514 8046
rect 96462 7970 96514 7982
rect 97246 8034 97298 8046
rect 97246 7970 97298 7982
rect 102398 8034 102450 8046
rect 102398 7970 102450 7982
rect 105086 8034 105138 8046
rect 105086 7970 105138 7982
rect 105758 8034 105810 8046
rect 105758 7970 105810 7982
rect 106206 8034 106258 8046
rect 106206 7970 106258 7982
rect 106654 8034 106706 8046
rect 106654 7970 106706 7982
rect 107998 8034 108050 8046
rect 112814 8034 112866 8046
rect 112242 7982 112254 8034
rect 112306 7982 112318 8034
rect 107998 7970 108050 7982
rect 112814 7970 112866 7982
rect 114158 8034 114210 8046
rect 114158 7970 114210 7982
rect 115166 8034 115218 8046
rect 115166 7970 115218 7982
rect 115726 8034 115778 8046
rect 115726 7970 115778 7982
rect 117854 8034 117906 8046
rect 117854 7970 117906 7982
rect 118302 8034 118354 8046
rect 118302 7970 118354 7982
rect 118862 8034 118914 8046
rect 121102 8034 121154 8046
rect 120194 7982 120206 8034
rect 120258 7982 120270 8034
rect 118862 7970 118914 7982
rect 121102 7970 121154 7982
rect 121550 8034 121602 8046
rect 121550 7970 121602 7982
rect 121998 8034 122050 8046
rect 121998 7970 122050 7982
rect 122558 8034 122610 8046
rect 122558 7970 122610 7982
rect 123006 8034 123058 8046
rect 123006 7970 123058 7982
rect 123790 8034 123842 8046
rect 123790 7970 123842 7982
rect 124350 8034 124402 8046
rect 124350 7970 124402 7982
rect 128830 8034 128882 8046
rect 128830 7970 128882 7982
rect 130622 8034 130674 8046
rect 130622 7970 130674 7982
rect 131070 8034 131122 8046
rect 131070 7970 131122 7982
rect 131406 8034 131458 8046
rect 131406 7970 131458 7982
rect 131966 8034 132018 8046
rect 131966 7970 132018 7982
rect 132974 8034 133026 8046
rect 132974 7970 133026 7982
rect 133646 8034 133698 8046
rect 133646 7970 133698 7982
rect 135102 8034 135154 8046
rect 135102 7970 135154 7982
rect 135438 8034 135490 8046
rect 135438 7970 135490 7982
rect 136670 8034 136722 8046
rect 136670 7970 136722 7982
rect 137566 8034 137618 8046
rect 137566 7970 137618 7982
rect 139694 8034 139746 8046
rect 139694 7970 139746 7982
rect 140142 8034 140194 8046
rect 140142 7970 140194 7982
rect 140926 8034 140978 8046
rect 140926 7970 140978 7982
rect 1344 7866 178640 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 81278 7866
rect 81330 7814 81382 7866
rect 81434 7814 81486 7866
rect 81538 7814 111998 7866
rect 112050 7814 112102 7866
rect 112154 7814 112206 7866
rect 112258 7814 142718 7866
rect 142770 7814 142822 7866
rect 142874 7814 142926 7866
rect 142978 7814 173438 7866
rect 173490 7814 173542 7866
rect 173594 7814 173646 7866
rect 173698 7814 178640 7866
rect 1344 7780 178640 7814
rect 31950 7698 32002 7710
rect 31950 7634 32002 7646
rect 37886 7698 37938 7710
rect 37886 7634 37938 7646
rect 39230 7698 39282 7710
rect 39230 7634 39282 7646
rect 47294 7698 47346 7710
rect 47294 7634 47346 7646
rect 55694 7698 55746 7710
rect 55694 7634 55746 7646
rect 61742 7698 61794 7710
rect 61742 7634 61794 7646
rect 62414 7698 62466 7710
rect 62414 7634 62466 7646
rect 73390 7698 73442 7710
rect 73390 7634 73442 7646
rect 75406 7698 75458 7710
rect 81678 7698 81730 7710
rect 80098 7646 80110 7698
rect 80162 7646 80174 7698
rect 75406 7634 75458 7646
rect 81678 7634 81730 7646
rect 90862 7698 90914 7710
rect 90862 7634 90914 7646
rect 91758 7698 91810 7710
rect 91758 7634 91810 7646
rect 93102 7698 93154 7710
rect 93102 7634 93154 7646
rect 93550 7698 93602 7710
rect 93550 7634 93602 7646
rect 93998 7698 94050 7710
rect 93998 7634 94050 7646
rect 94446 7698 94498 7710
rect 94446 7634 94498 7646
rect 94894 7698 94946 7710
rect 94894 7634 94946 7646
rect 97806 7698 97858 7710
rect 97806 7634 97858 7646
rect 98366 7698 98418 7710
rect 98366 7634 98418 7646
rect 99710 7698 99762 7710
rect 99710 7634 99762 7646
rect 100046 7698 100098 7710
rect 100046 7634 100098 7646
rect 100942 7698 100994 7710
rect 100942 7634 100994 7646
rect 101502 7698 101554 7710
rect 101502 7634 101554 7646
rect 102398 7698 102450 7710
rect 102398 7634 102450 7646
rect 103406 7698 103458 7710
rect 103406 7634 103458 7646
rect 103518 7698 103570 7710
rect 103518 7634 103570 7646
rect 104302 7698 104354 7710
rect 104302 7634 104354 7646
rect 105534 7698 105586 7710
rect 105534 7634 105586 7646
rect 106878 7698 106930 7710
rect 106878 7634 106930 7646
rect 107438 7698 107490 7710
rect 107438 7634 107490 7646
rect 109566 7698 109618 7710
rect 109566 7634 109618 7646
rect 109902 7698 109954 7710
rect 114382 7698 114434 7710
rect 112354 7646 112366 7698
rect 112418 7646 112430 7698
rect 109902 7634 109954 7646
rect 114382 7634 114434 7646
rect 114830 7698 114882 7710
rect 114830 7634 114882 7646
rect 115838 7698 115890 7710
rect 115838 7634 115890 7646
rect 120990 7698 121042 7710
rect 120990 7634 121042 7646
rect 123230 7698 123282 7710
rect 123230 7634 123282 7646
rect 124238 7698 124290 7710
rect 124238 7634 124290 7646
rect 129950 7698 130002 7710
rect 129950 7634 130002 7646
rect 130846 7698 130898 7710
rect 130846 7634 130898 7646
rect 131518 7698 131570 7710
rect 131518 7634 131570 7646
rect 132414 7698 132466 7710
rect 132414 7634 132466 7646
rect 134430 7698 134482 7710
rect 134430 7634 134482 7646
rect 137790 7698 137842 7710
rect 137790 7634 137842 7646
rect 138798 7698 138850 7710
rect 138798 7634 138850 7646
rect 32286 7586 32338 7598
rect 18946 7534 18958 7586
rect 19010 7534 19022 7586
rect 26450 7534 26462 7586
rect 26514 7534 26526 7586
rect 32286 7522 32338 7534
rect 39566 7586 39618 7598
rect 39566 7522 39618 7534
rect 42814 7586 42866 7598
rect 62862 7586 62914 7598
rect 73726 7586 73778 7598
rect 44146 7534 44158 7586
rect 44210 7534 44222 7586
rect 51090 7534 51102 7586
rect 51154 7534 51166 7586
rect 56018 7534 56030 7586
rect 56082 7583 56094 7586
rect 56242 7583 56254 7586
rect 56082 7537 56254 7583
rect 56082 7534 56094 7537
rect 56242 7534 56254 7537
rect 56306 7534 56318 7586
rect 69010 7534 69022 7586
rect 69074 7534 69086 7586
rect 42814 7522 42866 7534
rect 62862 7522 62914 7534
rect 73726 7522 73778 7534
rect 74286 7586 74338 7598
rect 78990 7586 79042 7598
rect 76514 7534 76526 7586
rect 76578 7534 76590 7586
rect 74286 7522 74338 7534
rect 78990 7522 79042 7534
rect 81566 7586 81618 7598
rect 95006 7586 95058 7598
rect 83906 7534 83918 7586
rect 83970 7534 83982 7586
rect 85026 7534 85038 7586
rect 85090 7534 85102 7586
rect 81566 7522 81618 7534
rect 95006 7522 95058 7534
rect 95230 7586 95282 7598
rect 95230 7522 95282 7534
rect 95678 7586 95730 7598
rect 95678 7522 95730 7534
rect 97358 7586 97410 7598
rect 104190 7586 104242 7598
rect 101826 7534 101838 7586
rect 101890 7534 101902 7586
rect 97358 7522 97410 7534
rect 104190 7522 104242 7534
rect 107998 7586 108050 7598
rect 107998 7522 108050 7534
rect 108110 7586 108162 7598
rect 108110 7522 108162 7534
rect 113150 7586 113202 7598
rect 113150 7522 113202 7534
rect 115950 7586 116002 7598
rect 115950 7522 116002 7534
rect 117630 7586 117682 7598
rect 117630 7522 117682 7534
rect 118190 7586 118242 7598
rect 118190 7522 118242 7534
rect 118414 7586 118466 7598
rect 118414 7522 118466 7534
rect 121438 7586 121490 7598
rect 121438 7522 121490 7534
rect 33518 7474 33570 7486
rect 37550 7474 37602 7486
rect 18274 7422 18286 7474
rect 18338 7422 18350 7474
rect 25666 7422 25678 7474
rect 25730 7422 25742 7474
rect 34178 7422 34190 7474
rect 34242 7422 34254 7474
rect 36082 7422 36094 7474
rect 36146 7422 36158 7474
rect 33518 7410 33570 7422
rect 37550 7410 37602 7422
rect 42478 7474 42530 7486
rect 46958 7474 47010 7486
rect 43362 7422 43374 7474
rect 43426 7422 43438 7474
rect 42478 7410 42530 7422
rect 46958 7410 47010 7422
rect 47854 7474 47906 7486
rect 55358 7474 55410 7486
rect 53890 7422 53902 7474
rect 53954 7422 53966 7474
rect 47854 7410 47906 7422
rect 55358 7410 55410 7422
rect 56366 7474 56418 7486
rect 62302 7474 62354 7486
rect 56690 7422 56702 7474
rect 56754 7422 56766 7474
rect 57810 7422 57822 7474
rect 57874 7422 57886 7474
rect 56366 7410 56418 7422
rect 62302 7410 62354 7422
rect 62526 7474 62578 7486
rect 62526 7410 62578 7422
rect 63422 7474 63474 7486
rect 63422 7410 63474 7422
rect 63646 7474 63698 7486
rect 63646 7410 63698 7422
rect 63870 7474 63922 7486
rect 75294 7474 75346 7486
rect 78542 7474 78594 7486
rect 89518 7474 89570 7486
rect 95454 7474 95506 7486
rect 66882 7422 66894 7474
rect 66946 7422 66958 7474
rect 71586 7422 71598 7474
rect 71650 7422 71662 7474
rect 74498 7422 74510 7474
rect 74562 7422 74574 7474
rect 76402 7422 76414 7474
rect 76466 7422 76478 7474
rect 82338 7422 82350 7474
rect 82402 7422 82414 7474
rect 84802 7422 84814 7474
rect 84866 7422 84878 7474
rect 86818 7422 86830 7474
rect 86882 7422 86894 7474
rect 89842 7422 89854 7474
rect 89906 7422 89918 7474
rect 63870 7410 63922 7422
rect 75294 7410 75346 7422
rect 78542 7410 78594 7422
rect 89518 7410 89570 7422
rect 95454 7410 95506 7422
rect 100494 7474 100546 7486
rect 100494 7410 100546 7422
rect 102734 7474 102786 7486
rect 102734 7410 102786 7422
rect 106430 7474 106482 7486
rect 106430 7410 106482 7422
rect 107774 7474 107826 7486
rect 107774 7410 107826 7422
rect 110798 7474 110850 7486
rect 110798 7410 110850 7422
rect 112030 7474 112082 7486
rect 115390 7474 115442 7486
rect 113362 7422 113374 7474
rect 113426 7422 113438 7474
rect 112030 7410 112082 7422
rect 115390 7410 115442 7422
rect 115614 7474 115666 7486
rect 115614 7410 115666 7422
rect 117294 7474 117346 7486
rect 117294 7410 117346 7422
rect 118750 7474 118802 7486
rect 130398 7474 130450 7486
rect 119634 7422 119646 7474
rect 119698 7422 119710 7474
rect 118750 7410 118802 7422
rect 130398 7410 130450 7422
rect 131966 7474 132018 7486
rect 131966 7410 132018 7422
rect 14926 7362 14978 7374
rect 14926 7298 14978 7310
rect 16382 7362 16434 7374
rect 21534 7362 21586 7374
rect 21074 7310 21086 7362
rect 21138 7310 21150 7362
rect 16382 7298 16434 7310
rect 21534 7298 21586 7310
rect 21982 7362 22034 7374
rect 21982 7298 22034 7310
rect 22430 7362 22482 7374
rect 22430 7298 22482 7310
rect 22878 7362 22930 7374
rect 22878 7298 22930 7310
rect 23438 7362 23490 7374
rect 23438 7298 23490 7310
rect 23886 7362 23938 7374
rect 23886 7298 23938 7310
rect 24222 7362 24274 7374
rect 29038 7362 29090 7374
rect 28578 7310 28590 7362
rect 28642 7310 28654 7362
rect 24222 7298 24274 7310
rect 29038 7298 29090 7310
rect 29598 7362 29650 7374
rect 29598 7298 29650 7310
rect 30046 7362 30098 7374
rect 30046 7298 30098 7310
rect 30606 7362 30658 7374
rect 30606 7298 30658 7310
rect 30942 7362 30994 7374
rect 30942 7298 30994 7310
rect 31502 7362 31554 7374
rect 31502 7298 31554 7310
rect 32846 7362 32898 7374
rect 32846 7298 32898 7310
rect 34638 7362 34690 7374
rect 34638 7298 34690 7310
rect 35310 7362 35362 7374
rect 35310 7298 35362 7310
rect 36654 7362 36706 7374
rect 36654 7298 36706 7310
rect 36990 7362 37042 7374
rect 36990 7298 37042 7310
rect 38782 7362 38834 7374
rect 38782 7298 38834 7310
rect 40462 7362 40514 7374
rect 40462 7298 40514 7310
rect 40910 7362 40962 7374
rect 40910 7298 40962 7310
rect 41582 7362 41634 7374
rect 41582 7298 41634 7310
rect 41918 7362 41970 7374
rect 48414 7362 48466 7374
rect 61406 7362 61458 7374
rect 46274 7310 46286 7362
rect 46338 7310 46350 7362
rect 58594 7310 58606 7362
rect 58658 7310 58670 7362
rect 60722 7310 60734 7362
rect 60786 7310 60798 7362
rect 41918 7298 41970 7310
rect 48414 7298 48466 7310
rect 61406 7298 61458 7310
rect 63534 7362 63586 7374
rect 63534 7298 63586 7310
rect 64654 7362 64706 7374
rect 87278 7362 87330 7374
rect 71698 7310 71710 7362
rect 71762 7310 71774 7362
rect 83122 7310 83134 7362
rect 83186 7310 83198 7362
rect 86482 7310 86494 7362
rect 86546 7310 86558 7362
rect 64654 7298 64706 7310
rect 87278 7298 87330 7310
rect 87726 7362 87778 7374
rect 87726 7298 87778 7310
rect 88510 7362 88562 7374
rect 88510 7298 88562 7310
rect 90414 7362 90466 7374
rect 90414 7298 90466 7310
rect 92094 7362 92146 7374
rect 92094 7298 92146 7310
rect 92766 7362 92818 7374
rect 92766 7298 92818 7310
rect 96126 7362 96178 7374
rect 96126 7298 96178 7310
rect 97246 7362 97298 7374
rect 97246 7298 97298 7310
rect 98702 7362 98754 7374
rect 98702 7298 98754 7310
rect 99150 7362 99202 7374
rect 99150 7298 99202 7310
rect 105086 7362 105138 7374
rect 105086 7298 105138 7310
rect 105982 7362 106034 7374
rect 105982 7298 106034 7310
rect 108558 7362 108610 7374
rect 108558 7298 108610 7310
rect 109006 7362 109058 7374
rect 109006 7298 109058 7310
rect 110350 7362 110402 7374
rect 110350 7298 110402 7310
rect 111246 7362 111298 7374
rect 111246 7298 111298 7310
rect 113934 7362 113986 7374
rect 113934 7298 113986 7310
rect 116398 7362 116450 7374
rect 116398 7298 116450 7310
rect 118638 7362 118690 7374
rect 120318 7362 120370 7374
rect 119410 7310 119422 7362
rect 119474 7310 119486 7362
rect 118638 7298 118690 7310
rect 120318 7298 120370 7310
rect 121998 7362 122050 7374
rect 121998 7298 122050 7310
rect 122446 7362 122498 7374
rect 122446 7298 122498 7310
rect 122894 7362 122946 7374
rect 122894 7298 122946 7310
rect 123790 7362 123842 7374
rect 123790 7298 123842 7310
rect 124686 7362 124738 7374
rect 124686 7298 124738 7310
rect 125022 7362 125074 7374
rect 125022 7298 125074 7310
rect 125470 7362 125522 7374
rect 125470 7298 125522 7310
rect 126142 7362 126194 7374
rect 126142 7298 126194 7310
rect 126478 7362 126530 7374
rect 126478 7298 126530 7310
rect 127934 7362 127986 7374
rect 127934 7298 127986 7310
rect 128382 7362 128434 7374
rect 128382 7298 128434 7310
rect 128942 7362 128994 7374
rect 128942 7298 128994 7310
rect 129502 7362 129554 7374
rect 129502 7298 129554 7310
rect 132750 7362 132802 7374
rect 132750 7298 132802 7310
rect 133198 7362 133250 7374
rect 133198 7298 133250 7310
rect 134094 7362 134146 7374
rect 134094 7298 134146 7310
rect 135214 7362 135266 7374
rect 135214 7298 135266 7310
rect 135662 7362 135714 7374
rect 135662 7298 135714 7310
rect 136110 7362 136162 7374
rect 136110 7298 136162 7310
rect 136894 7362 136946 7374
rect 136894 7298 136946 7310
rect 137342 7362 137394 7374
rect 137342 7298 137394 7310
rect 138238 7362 138290 7374
rect 138238 7298 138290 7310
rect 139134 7362 139186 7374
rect 139134 7298 139186 7310
rect 140030 7362 140082 7374
rect 140030 7298 140082 7310
rect 140478 7362 140530 7374
rect 140478 7298 140530 7310
rect 140926 7362 140978 7374
rect 140926 7298 140978 7310
rect 141598 7362 141650 7374
rect 141598 7298 141650 7310
rect 141934 7362 141986 7374
rect 141934 7298 141986 7310
rect 142718 7362 142770 7374
rect 142718 7298 142770 7310
rect 143054 7362 143106 7374
rect 143054 7298 143106 7310
rect 143614 7362 143666 7374
rect 143614 7298 143666 7310
rect 144846 7362 144898 7374
rect 144846 7298 144898 7310
rect 145406 7362 145458 7374
rect 145406 7298 145458 7310
rect 35758 7250 35810 7262
rect 35758 7186 35810 7198
rect 36094 7250 36146 7262
rect 36094 7186 36146 7198
rect 56702 7250 56754 7262
rect 75406 7250 75458 7262
rect 72370 7198 72382 7250
rect 72434 7198 72446 7250
rect 56702 7186 56754 7198
rect 75406 7186 75458 7198
rect 81678 7250 81730 7262
rect 81678 7186 81730 7198
rect 103294 7250 103346 7262
rect 109330 7198 109342 7250
rect 109394 7247 109406 7250
rect 110002 7247 110014 7250
rect 109394 7201 110014 7247
rect 109394 7198 109406 7201
rect 110002 7198 110014 7201
rect 110066 7198 110078 7250
rect 124450 7198 124462 7250
rect 124514 7247 124526 7250
rect 124674 7247 124686 7250
rect 124514 7201 124686 7247
rect 124514 7198 124526 7201
rect 124674 7198 124686 7201
rect 124738 7198 124750 7250
rect 132850 7198 132862 7250
rect 132914 7247 132926 7250
rect 133186 7247 133198 7250
rect 132914 7201 133198 7247
rect 132914 7198 132926 7201
rect 133186 7198 133198 7201
rect 133250 7198 133262 7250
rect 136770 7198 136782 7250
rect 136834 7247 136846 7250
rect 137778 7247 137790 7250
rect 136834 7201 137790 7247
rect 136834 7198 136846 7201
rect 137778 7198 137790 7201
rect 137842 7198 137854 7250
rect 103294 7186 103346 7198
rect 1344 7082 178640 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 96638 7082
rect 96690 7030 96742 7082
rect 96794 7030 96846 7082
rect 96898 7030 127358 7082
rect 127410 7030 127462 7082
rect 127514 7030 127566 7082
rect 127618 7030 158078 7082
rect 158130 7030 158182 7082
rect 158234 7030 158286 7082
rect 158338 7030 178640 7082
rect 1344 6996 178640 7030
rect 19630 6914 19682 6926
rect 19630 6850 19682 6862
rect 19966 6914 20018 6926
rect 19966 6850 20018 6862
rect 27470 6914 27522 6926
rect 27470 6850 27522 6862
rect 45950 6914 46002 6926
rect 45950 6850 46002 6862
rect 50430 6914 50482 6926
rect 50430 6850 50482 6862
rect 77758 6914 77810 6926
rect 77758 6850 77810 6862
rect 83134 6914 83186 6926
rect 83134 6850 83186 6862
rect 83470 6914 83522 6926
rect 135774 6914 135826 6926
rect 87490 6862 87502 6914
rect 87554 6911 87566 6914
rect 87714 6911 87726 6914
rect 87554 6865 87726 6911
rect 87554 6862 87566 6865
rect 87714 6862 87726 6865
rect 87778 6862 87790 6914
rect 91186 6862 91198 6914
rect 91250 6911 91262 6914
rect 91746 6911 91758 6914
rect 91250 6865 91758 6911
rect 91250 6862 91262 6865
rect 91746 6862 91758 6865
rect 91810 6862 91822 6914
rect 141586 6862 141598 6914
rect 141650 6911 141662 6914
rect 142146 6911 142158 6914
rect 141650 6865 142158 6911
rect 141650 6862 141662 6865
rect 142146 6862 142158 6865
rect 142210 6862 142222 6914
rect 143042 6862 143054 6914
rect 143106 6911 143118 6914
rect 143826 6911 143838 6914
rect 143106 6865 143838 6911
rect 143106 6862 143118 6865
rect 143826 6862 143838 6865
rect 143890 6862 143902 6914
rect 83470 6850 83522 6862
rect 135774 6850 135826 6862
rect 27806 6802 27858 6814
rect 76526 6802 76578 6814
rect 32050 6750 32062 6802
rect 32114 6750 32126 6802
rect 56354 6750 56366 6802
rect 56418 6750 56430 6802
rect 62962 6750 62974 6802
rect 63026 6750 63038 6802
rect 65090 6750 65102 6802
rect 65154 6750 65166 6802
rect 73826 6750 73838 6802
rect 73890 6750 73902 6802
rect 27806 6738 27858 6750
rect 76526 6738 76578 6750
rect 77534 6802 77586 6814
rect 87726 6802 87778 6814
rect 80658 6750 80670 6802
rect 80722 6750 80734 6802
rect 85810 6750 85822 6802
rect 85874 6750 85886 6802
rect 77534 6738 77586 6750
rect 87726 6738 87778 6750
rect 89742 6802 89794 6814
rect 89742 6738 89794 6750
rect 95118 6802 95170 6814
rect 95118 6738 95170 6750
rect 96686 6802 96738 6814
rect 101502 6802 101554 6814
rect 114382 6802 114434 6814
rect 119086 6802 119138 6814
rect 122894 6802 122946 6814
rect 97346 6750 97358 6802
rect 97410 6750 97422 6802
rect 102722 6750 102734 6802
rect 102786 6750 102798 6802
rect 105858 6750 105870 6802
rect 105922 6750 105934 6802
rect 109330 6750 109342 6802
rect 109394 6750 109406 6802
rect 115490 6750 115502 6802
rect 115554 6750 115566 6802
rect 120194 6750 120206 6802
rect 120258 6750 120270 6802
rect 96686 6738 96738 6750
rect 101502 6738 101554 6750
rect 114382 6738 114434 6750
rect 119086 6738 119138 6750
rect 122894 6738 122946 6750
rect 35982 6690 36034 6702
rect 20626 6638 20638 6690
rect 20690 6638 20702 6690
rect 24098 6638 24110 6690
rect 24162 6638 24174 6690
rect 25890 6638 25902 6690
rect 25954 6638 25966 6690
rect 34850 6638 34862 6690
rect 34914 6638 34926 6690
rect 35982 6626 36034 6638
rect 36430 6690 36482 6702
rect 36430 6626 36482 6638
rect 37438 6690 37490 6702
rect 37438 6626 37490 6638
rect 37774 6690 37826 6702
rect 42366 6690 42418 6702
rect 43374 6690 43426 6702
rect 45614 6690 45666 6702
rect 50766 6690 50818 6702
rect 57150 6690 57202 6702
rect 65886 6690 65938 6702
rect 38882 6638 38894 6690
rect 38946 6638 38958 6690
rect 42914 6638 42926 6690
rect 42978 6638 42990 6690
rect 44594 6638 44606 6690
rect 44658 6638 44670 6690
rect 46722 6638 46734 6690
rect 46786 6638 46798 6690
rect 49746 6638 49758 6690
rect 49810 6638 49822 6690
rect 51426 6638 51438 6690
rect 51490 6638 51502 6690
rect 53442 6638 53454 6690
rect 53506 6638 53518 6690
rect 54226 6638 54238 6690
rect 54290 6638 54302 6690
rect 62178 6638 62190 6690
rect 62242 6638 62254 6690
rect 37774 6626 37826 6638
rect 42366 6626 42418 6638
rect 43374 6626 43426 6638
rect 45614 6626 45666 6638
rect 50766 6626 50818 6638
rect 57150 6626 57202 6638
rect 65886 6626 65938 6638
rect 66110 6690 66162 6702
rect 66110 6626 66162 6638
rect 66334 6690 66386 6702
rect 66334 6626 66386 6638
rect 66558 6690 66610 6702
rect 66558 6626 66610 6638
rect 68574 6690 68626 6702
rect 79662 6690 79714 6702
rect 82126 6690 82178 6702
rect 69346 6638 69358 6690
rect 69410 6638 69422 6690
rect 77298 6638 77310 6690
rect 77362 6638 77374 6690
rect 80770 6638 80782 6690
rect 80834 6638 80846 6690
rect 68574 6626 68626 6638
rect 79662 6626 79714 6638
rect 82126 6626 82178 6638
rect 82910 6690 82962 6702
rect 87278 6690 87330 6702
rect 85250 6638 85262 6690
rect 85314 6638 85326 6690
rect 82910 6626 82962 6638
rect 87278 6626 87330 6638
rect 89294 6690 89346 6702
rect 89294 6626 89346 6638
rect 91534 6690 91586 6702
rect 91534 6626 91586 6638
rect 91982 6690 92034 6702
rect 91982 6626 92034 6638
rect 92318 6690 92370 6702
rect 92318 6626 92370 6638
rect 93102 6690 93154 6702
rect 93102 6626 93154 6638
rect 93774 6690 93826 6702
rect 93774 6626 93826 6638
rect 95678 6690 95730 6702
rect 95678 6626 95730 6638
rect 95902 6690 95954 6702
rect 95902 6626 95954 6638
rect 96238 6690 96290 6702
rect 99486 6690 99538 6702
rect 97458 6638 97470 6690
rect 97522 6638 97534 6690
rect 97682 6638 97694 6690
rect 97746 6638 97758 6690
rect 96238 6626 96290 6638
rect 99486 6626 99538 6638
rect 99934 6690 99986 6702
rect 99934 6626 99986 6638
rect 101054 6690 101106 6702
rect 103966 6690 104018 6702
rect 102610 6638 102622 6690
rect 102674 6638 102686 6690
rect 101054 6626 101106 6638
rect 103966 6626 104018 6638
rect 104190 6690 104242 6702
rect 110238 6690 110290 6702
rect 105074 6638 105086 6690
rect 105138 6638 105150 6690
rect 106754 6638 106766 6690
rect 106818 6638 106830 6690
rect 104190 6626 104242 6638
rect 110238 6626 110290 6638
rect 111134 6690 111186 6702
rect 111134 6626 111186 6638
rect 112142 6690 112194 6702
rect 112142 6626 112194 6638
rect 113934 6690 113986 6702
rect 113934 6626 113986 6638
rect 117406 6690 117458 6702
rect 117406 6626 117458 6638
rect 119310 6690 119362 6702
rect 122446 6690 122498 6702
rect 120418 6638 120430 6690
rect 120482 6638 120494 6690
rect 119310 6626 119362 6638
rect 122446 6626 122498 6638
rect 123902 6690 123954 6702
rect 123902 6626 123954 6638
rect 126926 6690 126978 6702
rect 126926 6626 126978 6638
rect 128046 6690 128098 6702
rect 128046 6626 128098 6638
rect 128606 6690 128658 6702
rect 128606 6626 128658 6638
rect 128942 6690 128994 6702
rect 130622 6690 130674 6702
rect 132302 6690 132354 6702
rect 130050 6638 130062 6690
rect 130114 6638 130126 6690
rect 130946 6638 130958 6690
rect 131010 6638 131022 6690
rect 128942 6626 128994 6638
rect 130622 6626 130674 6638
rect 132302 6626 132354 6638
rect 135886 6690 135938 6702
rect 135886 6626 135938 6638
rect 141262 6690 141314 6702
rect 141262 6626 141314 6638
rect 143950 6690 144002 6702
rect 143950 6626 144002 6638
rect 14590 6578 14642 6590
rect 14590 6514 14642 6526
rect 18734 6578 18786 6590
rect 21534 6578 21586 6590
rect 20738 6526 20750 6578
rect 20802 6526 20814 6578
rect 18734 6514 18786 6526
rect 21534 6514 21586 6526
rect 22654 6578 22706 6590
rect 29598 6578 29650 6590
rect 24322 6526 24334 6578
rect 24386 6526 24398 6578
rect 28130 6526 28142 6578
rect 28194 6526 28206 6578
rect 28578 6526 28590 6578
rect 28642 6526 28654 6578
rect 22654 6514 22706 6526
rect 29598 6514 29650 6526
rect 29934 6578 29986 6590
rect 29934 6514 29986 6526
rect 30494 6578 30546 6590
rect 35758 6578 35810 6590
rect 34178 6526 34190 6578
rect 34242 6526 34254 6578
rect 30494 6514 30546 6526
rect 35758 6514 35810 6526
rect 36206 6578 36258 6590
rect 36206 6514 36258 6526
rect 38110 6578 38162 6590
rect 38110 6514 38162 6526
rect 39678 6578 39730 6590
rect 39678 6514 39730 6526
rect 40014 6578 40066 6590
rect 40014 6514 40066 6526
rect 40574 6578 40626 6590
rect 40574 6514 40626 6526
rect 40910 6578 40962 6590
rect 40910 6514 40962 6526
rect 41806 6578 41858 6590
rect 41806 6514 41858 6526
rect 42590 6578 42642 6590
rect 44382 6578 44434 6590
rect 47742 6578 47794 6590
rect 42802 6526 42814 6578
rect 42866 6526 42878 6578
rect 46498 6526 46510 6578
rect 46562 6526 46574 6578
rect 42590 6514 42642 6526
rect 44382 6514 44434 6526
rect 47742 6514 47794 6526
rect 48078 6578 48130 6590
rect 48078 6514 48130 6526
rect 48638 6578 48690 6590
rect 48638 6514 48690 6526
rect 48974 6578 49026 6590
rect 57710 6578 57762 6590
rect 49634 6526 49646 6578
rect 49698 6526 49710 6578
rect 52322 6526 52334 6578
rect 52386 6526 52398 6578
rect 48974 6514 49026 6526
rect 57710 6514 57762 6526
rect 58046 6578 58098 6590
rect 58046 6514 58098 6526
rect 59390 6578 59442 6590
rect 59390 6514 59442 6526
rect 60622 6578 60674 6590
rect 60622 6514 60674 6526
rect 67678 6578 67730 6590
rect 67678 6514 67730 6526
rect 68126 6578 68178 6590
rect 68126 6514 68178 6526
rect 75518 6578 75570 6590
rect 75518 6514 75570 6526
rect 78430 6578 78482 6590
rect 78430 6514 78482 6526
rect 78766 6578 78818 6590
rect 78766 6514 78818 6526
rect 79774 6578 79826 6590
rect 79774 6514 79826 6526
rect 81454 6578 81506 6590
rect 81454 6514 81506 6526
rect 82238 6578 82290 6590
rect 82238 6514 82290 6526
rect 84478 6578 84530 6590
rect 84478 6514 84530 6526
rect 85822 6578 85874 6590
rect 85822 6514 85874 6526
rect 86830 6578 86882 6590
rect 86830 6514 86882 6526
rect 97246 6578 97298 6590
rect 97246 6514 97298 6526
rect 98590 6578 98642 6590
rect 98590 6514 98642 6526
rect 99038 6578 99090 6590
rect 99038 6514 99090 6526
rect 103070 6578 103122 6590
rect 109118 6578 109170 6590
rect 104514 6526 104526 6578
rect 104578 6526 104590 6578
rect 105634 6526 105646 6578
rect 105698 6526 105710 6578
rect 106642 6526 106654 6578
rect 106706 6526 106718 6578
rect 103070 6514 103122 6526
rect 109118 6514 109170 6526
rect 113038 6578 113090 6590
rect 115950 6578 116002 6590
rect 115714 6526 115726 6578
rect 115778 6526 115790 6578
rect 113038 6514 113090 6526
rect 115950 6514 116002 6526
rect 116062 6578 116114 6590
rect 116062 6514 116114 6526
rect 117854 6578 117906 6590
rect 117854 6514 117906 6526
rect 121102 6578 121154 6590
rect 121102 6514 121154 6526
rect 129726 6578 129778 6590
rect 129726 6514 129778 6526
rect 136670 6578 136722 6590
rect 136670 6514 136722 6526
rect 139134 6578 139186 6590
rect 139134 6514 139186 6526
rect 14142 6466 14194 6478
rect 14142 6402 14194 6414
rect 14926 6466 14978 6478
rect 14926 6402 14978 6414
rect 15486 6466 15538 6478
rect 15486 6402 15538 6414
rect 15822 6466 15874 6478
rect 15822 6402 15874 6414
rect 16382 6466 16434 6478
rect 16382 6402 16434 6414
rect 16942 6466 16994 6478
rect 16942 6402 16994 6414
rect 17390 6466 17442 6478
rect 17390 6402 17442 6414
rect 17726 6466 17778 6478
rect 17726 6402 17778 6414
rect 18174 6466 18226 6478
rect 18174 6402 18226 6414
rect 18846 6466 18898 6478
rect 18846 6402 18898 6414
rect 19070 6466 19122 6478
rect 19070 6402 19122 6414
rect 22206 6466 22258 6478
rect 22206 6402 22258 6414
rect 23214 6466 23266 6478
rect 23214 6402 23266 6414
rect 24782 6466 24834 6478
rect 24782 6402 24834 6414
rect 25342 6466 25394 6478
rect 25342 6402 25394 6414
rect 26126 6466 26178 6478
rect 26126 6402 26178 6414
rect 26910 6466 26962 6478
rect 26910 6402 26962 6414
rect 31054 6466 31106 6478
rect 31054 6402 31106 6414
rect 31614 6466 31666 6478
rect 31614 6402 31666 6414
rect 36878 6466 36930 6478
rect 36878 6402 36930 6414
rect 37774 6466 37826 6478
rect 37774 6402 37826 6414
rect 39118 6466 39170 6478
rect 39118 6402 39170 6414
rect 41470 6466 41522 6478
rect 41470 6402 41522 6414
rect 43822 6466 43874 6478
rect 43822 6402 43874 6414
rect 58830 6466 58882 6478
rect 58830 6402 58882 6414
rect 59726 6466 59778 6478
rect 59726 6402 59778 6414
rect 60398 6466 60450 6478
rect 60398 6402 60450 6414
rect 60510 6466 60562 6478
rect 60510 6402 60562 6414
rect 61742 6466 61794 6478
rect 67902 6466 67954 6478
rect 66994 6414 67006 6466
rect 67058 6414 67070 6466
rect 61742 6402 61794 6414
rect 67902 6402 67954 6414
rect 68238 6466 68290 6478
rect 68238 6402 68290 6414
rect 75182 6466 75234 6478
rect 75182 6402 75234 6414
rect 76414 6466 76466 6478
rect 76414 6402 76466 6414
rect 77422 6466 77474 6478
rect 77422 6402 77474 6414
rect 79998 6466 80050 6478
rect 79998 6402 80050 6414
rect 82462 6466 82514 6478
rect 82462 6402 82514 6414
rect 84142 6466 84194 6478
rect 84142 6402 84194 6414
rect 85486 6466 85538 6478
rect 85486 6402 85538 6414
rect 85710 6466 85762 6478
rect 85710 6402 85762 6414
rect 86494 6466 86546 6478
rect 86494 6402 86546 6414
rect 88398 6466 88450 6478
rect 88398 6402 88450 6414
rect 90078 6466 90130 6478
rect 90078 6402 90130 6414
rect 90526 6466 90578 6478
rect 90526 6402 90578 6414
rect 90974 6466 91026 6478
rect 90974 6402 91026 6414
rect 94446 6466 94498 6478
rect 94446 6402 94498 6414
rect 95902 6466 95954 6478
rect 95902 6402 95954 6414
rect 98254 6466 98306 6478
rect 98254 6402 98306 6414
rect 100382 6466 100434 6478
rect 100382 6402 100434 6414
rect 109342 6466 109394 6478
rect 109342 6402 109394 6414
rect 110574 6466 110626 6478
rect 110574 6402 110626 6414
rect 111246 6466 111298 6478
rect 111246 6402 111298 6414
rect 111694 6466 111746 6478
rect 111694 6402 111746 6414
rect 112590 6466 112642 6478
rect 112590 6402 112642 6414
rect 113486 6466 113538 6478
rect 113486 6402 113538 6414
rect 114830 6466 114882 6478
rect 114830 6402 114882 6414
rect 116286 6466 116338 6478
rect 116286 6402 116338 6414
rect 117070 6466 117122 6478
rect 121550 6466 121602 6478
rect 118738 6414 118750 6466
rect 118802 6414 118814 6466
rect 117070 6402 117122 6414
rect 121550 6402 121602 6414
rect 121998 6466 122050 6478
rect 121998 6402 122050 6414
rect 123454 6466 123506 6478
rect 123454 6402 123506 6414
rect 124238 6466 124290 6478
rect 124238 6402 124290 6414
rect 124910 6466 124962 6478
rect 124910 6402 124962 6414
rect 125358 6466 125410 6478
rect 125358 6402 125410 6414
rect 125806 6466 125858 6478
rect 125806 6402 125858 6414
rect 126478 6466 126530 6478
rect 126478 6402 126530 6414
rect 127374 6466 127426 6478
rect 127374 6402 127426 6414
rect 129838 6466 129890 6478
rect 129838 6402 129890 6414
rect 130734 6466 130786 6478
rect 130734 6402 130786 6414
rect 131630 6466 131682 6478
rect 131630 6402 131682 6414
rect 133310 6466 133362 6478
rect 133310 6402 133362 6414
rect 133870 6466 133922 6478
rect 133870 6402 133922 6414
rect 134318 6466 134370 6478
rect 134318 6402 134370 6414
rect 134990 6466 135042 6478
rect 134990 6402 135042 6414
rect 135998 6466 136050 6478
rect 135998 6402 136050 6414
rect 137230 6466 137282 6478
rect 137230 6402 137282 6414
rect 137678 6466 137730 6478
rect 137678 6402 137730 6414
rect 138126 6466 138178 6478
rect 138126 6402 138178 6414
rect 138686 6466 138738 6478
rect 138686 6402 138738 6414
rect 139582 6466 139634 6478
rect 139582 6402 139634 6414
rect 139918 6466 139970 6478
rect 139918 6402 139970 6414
rect 140926 6466 140978 6478
rect 140926 6402 140978 6414
rect 141710 6466 141762 6478
rect 141710 6402 141762 6414
rect 142270 6466 142322 6478
rect 142270 6402 142322 6414
rect 142606 6466 142658 6478
rect 142606 6402 142658 6414
rect 143054 6466 143106 6478
rect 143054 6402 143106 6414
rect 143502 6466 143554 6478
rect 143502 6402 143554 6414
rect 144510 6466 144562 6478
rect 144510 6402 144562 6414
rect 145070 6466 145122 6478
rect 145070 6402 145122 6414
rect 145742 6466 145794 6478
rect 145742 6402 145794 6414
rect 146302 6466 146354 6478
rect 146302 6402 146354 6414
rect 146638 6466 146690 6478
rect 146638 6402 146690 6414
rect 147086 6466 147138 6478
rect 147086 6402 147138 6414
rect 147646 6466 147698 6478
rect 147646 6402 147698 6414
rect 148766 6466 148818 6478
rect 148766 6402 148818 6414
rect 1344 6298 178640 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 81278 6298
rect 81330 6246 81382 6298
rect 81434 6246 81486 6298
rect 81538 6246 111998 6298
rect 112050 6246 112102 6298
rect 112154 6246 112206 6298
rect 112258 6246 142718 6298
rect 142770 6246 142822 6298
rect 142874 6246 142926 6298
rect 142978 6246 173438 6298
rect 173490 6246 173542 6298
rect 173594 6246 173646 6298
rect 173698 6246 178640 6298
rect 1344 6212 178640 6246
rect 15262 6130 15314 6142
rect 15262 6066 15314 6078
rect 16046 6130 16098 6142
rect 16046 6066 16098 6078
rect 16718 6130 16770 6142
rect 16718 6066 16770 6078
rect 16942 6130 16994 6142
rect 16942 6066 16994 6078
rect 22766 6130 22818 6142
rect 22766 6066 22818 6078
rect 23550 6130 23602 6142
rect 23550 6066 23602 6078
rect 24446 6130 24498 6142
rect 24446 6066 24498 6078
rect 24894 6130 24946 6142
rect 24894 6066 24946 6078
rect 29150 6130 29202 6142
rect 29150 6066 29202 6078
rect 32846 6130 32898 6142
rect 32846 6066 32898 6078
rect 34974 6130 35026 6142
rect 34974 6066 35026 6078
rect 39342 6130 39394 6142
rect 39342 6066 39394 6078
rect 41918 6130 41970 6142
rect 41918 6066 41970 6078
rect 46062 6130 46114 6142
rect 46062 6066 46114 6078
rect 46846 6130 46898 6142
rect 46846 6066 46898 6078
rect 47742 6130 47794 6142
rect 47742 6066 47794 6078
rect 56590 6130 56642 6142
rect 56590 6066 56642 6078
rect 59390 6130 59442 6142
rect 59390 6066 59442 6078
rect 61630 6130 61682 6142
rect 65550 6130 65602 6142
rect 62850 6078 62862 6130
rect 62914 6078 62926 6130
rect 61630 6066 61682 6078
rect 65550 6066 65602 6078
rect 66558 6130 66610 6142
rect 66558 6066 66610 6078
rect 67678 6130 67730 6142
rect 67678 6066 67730 6078
rect 67790 6130 67842 6142
rect 67790 6066 67842 6078
rect 69470 6130 69522 6142
rect 69470 6066 69522 6078
rect 74734 6130 74786 6142
rect 74734 6066 74786 6078
rect 77758 6130 77810 6142
rect 77758 6066 77810 6078
rect 79886 6130 79938 6142
rect 79886 6066 79938 6078
rect 81454 6130 81506 6142
rect 81454 6066 81506 6078
rect 81678 6130 81730 6142
rect 81678 6066 81730 6078
rect 82350 6130 82402 6142
rect 82350 6066 82402 6078
rect 82574 6130 82626 6142
rect 82574 6066 82626 6078
rect 89182 6130 89234 6142
rect 89182 6066 89234 6078
rect 90750 6130 90802 6142
rect 90750 6066 90802 6078
rect 93102 6130 93154 6142
rect 93102 6066 93154 6078
rect 93662 6130 93714 6142
rect 93662 6066 93714 6078
rect 95006 6130 95058 6142
rect 99262 6130 99314 6142
rect 96114 6078 96126 6130
rect 96178 6078 96190 6130
rect 95006 6066 95058 6078
rect 99262 6066 99314 6078
rect 100718 6130 100770 6142
rect 103070 6130 103122 6142
rect 101714 6078 101726 6130
rect 101778 6078 101790 6130
rect 100718 6066 100770 6078
rect 103070 6066 103122 6078
rect 114046 6130 114098 6142
rect 114046 6066 114098 6078
rect 114382 6130 114434 6142
rect 114382 6066 114434 6078
rect 116062 6130 116114 6142
rect 116062 6066 116114 6078
rect 116958 6130 117010 6142
rect 116958 6066 117010 6078
rect 127262 6130 127314 6142
rect 127262 6066 127314 6078
rect 128046 6130 128098 6142
rect 128046 6066 128098 6078
rect 133870 6130 133922 6142
rect 133870 6066 133922 6078
rect 134654 6130 134706 6142
rect 134654 6066 134706 6078
rect 136222 6130 136274 6142
rect 136222 6066 136274 6078
rect 137006 6130 137058 6142
rect 137006 6066 137058 6078
rect 139918 6130 139970 6142
rect 139918 6066 139970 6078
rect 140814 6130 140866 6142
rect 140814 6066 140866 6078
rect 142494 6130 142546 6142
rect 142494 6066 142546 6078
rect 8430 6018 8482 6030
rect 8430 5954 8482 5966
rect 13470 6018 13522 6030
rect 13470 5954 13522 5966
rect 14366 6018 14418 6030
rect 14366 5954 14418 5966
rect 14926 6018 14978 6030
rect 14926 5954 14978 5966
rect 15038 6018 15090 6030
rect 20302 6018 20354 6030
rect 18386 5966 18398 6018
rect 18450 5966 18462 6018
rect 18946 5966 18958 6018
rect 19010 5966 19022 6018
rect 15038 5954 15090 5966
rect 20302 5954 20354 5966
rect 21534 6018 21586 6030
rect 34190 6018 34242 6030
rect 39230 6018 39282 6030
rect 26450 5966 26462 6018
rect 26514 5966 26526 6018
rect 37762 5966 37774 6018
rect 37826 5966 37838 6018
rect 21534 5954 21586 5966
rect 34190 5954 34242 5966
rect 39230 5954 39282 5966
rect 40462 6018 40514 6030
rect 40462 5954 40514 5966
rect 40798 6018 40850 6030
rect 42702 6018 42754 6030
rect 42466 5966 42478 6018
rect 42530 5966 42542 6018
rect 40798 5954 40850 5966
rect 42702 5954 42754 5966
rect 44158 6018 44210 6030
rect 44158 5954 44210 5966
rect 44606 6018 44658 6030
rect 44606 5954 44658 5966
rect 44830 6018 44882 6030
rect 44830 5954 44882 5966
rect 47630 6018 47682 6030
rect 47630 5954 47682 5966
rect 48862 6018 48914 6030
rect 57486 6018 57538 6030
rect 52210 5966 52222 6018
rect 52274 5966 52286 6018
rect 55682 5966 55694 6018
rect 55746 5966 55758 6018
rect 48862 5954 48914 5966
rect 57486 5954 57538 5966
rect 57710 6018 57762 6030
rect 57710 5954 57762 5966
rect 58046 6018 58098 6030
rect 58046 5954 58098 5966
rect 60734 6018 60786 6030
rect 60734 5954 60786 5966
rect 61294 6018 61346 6030
rect 61294 5954 61346 5966
rect 61518 6018 61570 6030
rect 61518 5954 61570 5966
rect 61854 6018 61906 6030
rect 61854 5954 61906 5966
rect 63422 6018 63474 6030
rect 63422 5954 63474 5966
rect 63646 6018 63698 6030
rect 63646 5954 63698 5966
rect 64318 6018 64370 6030
rect 64318 5954 64370 5966
rect 64654 6018 64706 6030
rect 64654 5954 64706 5966
rect 66110 6018 66162 6030
rect 66110 5954 66162 5966
rect 66334 6018 66386 6030
rect 66334 5954 66386 5966
rect 67230 6018 67282 6030
rect 67230 5954 67282 5966
rect 69358 6018 69410 6030
rect 69358 5954 69410 5966
rect 74062 6018 74114 6030
rect 74062 5954 74114 5966
rect 75182 6018 75234 6030
rect 75182 5954 75234 5966
rect 77646 6018 77698 6030
rect 77646 5954 77698 5966
rect 79102 6018 79154 6030
rect 79102 5954 79154 5966
rect 80446 6018 80498 6030
rect 80446 5954 80498 5966
rect 81342 6018 81394 6030
rect 81342 5954 81394 5966
rect 84030 6018 84082 6030
rect 84030 5954 84082 5966
rect 86046 6018 86098 6030
rect 86046 5954 86098 5966
rect 87838 6018 87890 6030
rect 87838 5954 87890 5966
rect 88174 6018 88226 6030
rect 88174 5954 88226 5966
rect 90414 6018 90466 6030
rect 90414 5954 90466 5966
rect 91646 6018 91698 6030
rect 91646 5954 91698 5966
rect 91870 6018 91922 6030
rect 91870 5954 91922 5966
rect 92542 6018 92594 6030
rect 92542 5954 92594 5966
rect 92654 6018 92706 6030
rect 92654 5954 92706 5966
rect 95566 6018 95618 6030
rect 99822 6018 99874 6030
rect 96226 5966 96238 6018
rect 96290 5966 96302 6018
rect 95566 5954 95618 5966
rect 99822 5954 99874 5966
rect 100158 6018 100210 6030
rect 102958 6018 103010 6030
rect 101826 5966 101838 6018
rect 101890 5966 101902 6018
rect 100158 5954 100210 5966
rect 102958 5954 103010 5966
rect 104078 6018 104130 6030
rect 104078 5954 104130 5966
rect 104414 6018 104466 6030
rect 104414 5954 104466 5966
rect 106878 6018 106930 6030
rect 106878 5954 106930 5966
rect 107102 6018 107154 6030
rect 107102 5954 107154 5966
rect 107998 6018 108050 6030
rect 107998 5954 108050 5966
rect 108334 6018 108386 6030
rect 108334 5954 108386 5966
rect 115278 6018 115330 6030
rect 115278 5954 115330 5966
rect 115614 6018 115666 6030
rect 115614 5954 115666 5966
rect 117630 6018 117682 6030
rect 117630 5954 117682 5966
rect 121214 6018 121266 6030
rect 121214 5954 121266 5966
rect 123118 6018 123170 6030
rect 123118 5954 123170 5966
rect 123790 6018 123842 6030
rect 123790 5954 123842 5966
rect 124910 6018 124962 6030
rect 124910 5954 124962 5966
rect 129054 6018 129106 6030
rect 129054 5954 129106 5966
rect 130846 6018 130898 6030
rect 130846 5954 130898 5966
rect 131182 6018 131234 6030
rect 131182 5954 131234 5966
rect 131742 6018 131794 6030
rect 131742 5954 131794 5966
rect 132638 6018 132690 6030
rect 132638 5954 132690 5966
rect 132974 6018 133026 6030
rect 132974 5954 133026 5966
rect 133758 6018 133810 6030
rect 133758 5954 133810 5966
rect 134542 6018 134594 6030
rect 134542 5954 134594 5966
rect 135774 6018 135826 6030
rect 135774 5954 135826 5966
rect 138350 6018 138402 6030
rect 138350 5954 138402 5966
rect 140702 6018 140754 6030
rect 140702 5954 140754 5966
rect 141710 6018 141762 6030
rect 141710 5954 141762 5966
rect 142382 6018 142434 6030
rect 142382 5954 142434 5966
rect 143390 6018 143442 6030
rect 143390 5954 143442 5966
rect 145294 6018 145346 6030
rect 145294 5954 145346 5966
rect 146750 6018 146802 6030
rect 146750 5954 146802 5966
rect 14030 5906 14082 5918
rect 8642 5854 8654 5906
rect 8706 5854 8718 5906
rect 13234 5854 13246 5906
rect 13298 5854 13310 5906
rect 14030 5842 14082 5854
rect 15710 5906 15762 5918
rect 15710 5842 15762 5854
rect 16606 5906 16658 5918
rect 16606 5842 16658 5854
rect 20638 5906 20690 5918
rect 20638 5842 20690 5854
rect 21198 5906 21250 5918
rect 21198 5842 21250 5854
rect 22430 5906 22482 5918
rect 22430 5842 22482 5854
rect 24110 5906 24162 5918
rect 33854 5906 33906 5918
rect 25666 5854 25678 5906
rect 25730 5854 25742 5906
rect 30930 5854 30942 5906
rect 30994 5854 31006 5906
rect 32610 5854 32622 5906
rect 32674 5854 32686 5906
rect 24110 5842 24162 5854
rect 33854 5842 33906 5854
rect 34750 5906 34802 5918
rect 39454 5906 39506 5918
rect 38546 5854 38558 5906
rect 38610 5854 38622 5906
rect 34750 5842 34802 5854
rect 39454 5842 39506 5854
rect 42366 5906 42418 5918
rect 45278 5906 45330 5918
rect 47406 5906 47458 5918
rect 42914 5854 42926 5906
rect 42978 5854 42990 5906
rect 46610 5854 46622 5906
rect 46674 5854 46686 5906
rect 42366 5842 42418 5854
rect 45278 5842 45330 5854
rect 47406 5842 47458 5854
rect 47966 5906 48018 5918
rect 56254 5906 56306 5918
rect 49970 5854 49982 5906
rect 50034 5854 50046 5906
rect 55458 5854 55470 5906
rect 55522 5854 55534 5906
rect 47966 5842 48018 5854
rect 56254 5842 56306 5854
rect 58942 5906 58994 5918
rect 58942 5842 58994 5854
rect 59614 5906 59666 5918
rect 59614 5842 59666 5854
rect 60398 5906 60450 5918
rect 60398 5842 60450 5854
rect 62526 5906 62578 5918
rect 62526 5842 62578 5854
rect 66782 5906 66834 5918
rect 66782 5842 66834 5854
rect 67454 5906 67506 5918
rect 67454 5842 67506 5854
rect 67566 5906 67618 5918
rect 68798 5906 68850 5918
rect 68450 5854 68462 5906
rect 68514 5854 68526 5906
rect 67566 5842 67618 5854
rect 68798 5842 68850 5854
rect 69134 5906 69186 5918
rect 69134 5842 69186 5854
rect 70030 5906 70082 5918
rect 72606 5906 72658 5918
rect 73614 5906 73666 5918
rect 70242 5854 70254 5906
rect 70306 5854 70318 5906
rect 71922 5854 71934 5906
rect 71986 5854 71998 5906
rect 73378 5854 73390 5906
rect 73442 5854 73454 5906
rect 70030 5842 70082 5854
rect 72606 5842 72658 5854
rect 73614 5842 73666 5854
rect 73950 5906 74002 5918
rect 73950 5842 74002 5854
rect 74398 5906 74450 5918
rect 77982 5906 78034 5918
rect 75394 5854 75406 5906
rect 75458 5854 75470 5906
rect 76514 5854 76526 5906
rect 76578 5854 76590 5906
rect 74398 5842 74450 5854
rect 77982 5842 78034 5854
rect 78094 5906 78146 5918
rect 80334 5906 80386 5918
rect 78866 5854 78878 5906
rect 78930 5854 78942 5906
rect 78094 5842 78146 5854
rect 80334 5842 80386 5854
rect 80670 5906 80722 5918
rect 82686 5906 82738 5918
rect 89966 5906 90018 5918
rect 82114 5854 82126 5906
rect 82178 5854 82190 5906
rect 83458 5854 83470 5906
rect 83522 5854 83534 5906
rect 85474 5854 85486 5906
rect 85538 5854 85550 5906
rect 89730 5854 89742 5906
rect 89794 5854 89806 5906
rect 80670 5842 80722 5854
rect 82686 5842 82738 5854
rect 89966 5842 90018 5854
rect 90078 5906 90130 5918
rect 90078 5842 90130 5854
rect 90750 5906 90802 5918
rect 90750 5842 90802 5854
rect 94670 5906 94722 5918
rect 97470 5906 97522 5918
rect 98926 5906 98978 5918
rect 102062 5906 102114 5918
rect 107438 5906 107490 5918
rect 113150 5906 113202 5918
rect 96450 5854 96462 5906
rect 96514 5854 96526 5906
rect 98130 5854 98142 5906
rect 98194 5854 98206 5906
rect 101266 5854 101278 5906
rect 101330 5854 101342 5906
rect 105634 5854 105646 5906
rect 105698 5854 105710 5906
rect 109218 5854 109230 5906
rect 109282 5854 109294 5906
rect 94670 5842 94722 5854
rect 97470 5842 97522 5854
rect 98926 5842 98978 5854
rect 102062 5842 102114 5854
rect 107438 5842 107490 5854
rect 113150 5842 113202 5854
rect 113374 5906 113426 5918
rect 113374 5842 113426 5854
rect 118414 5906 118466 5918
rect 118414 5842 118466 5854
rect 119758 5906 119810 5918
rect 119758 5842 119810 5854
rect 119870 5906 119922 5918
rect 128270 5906 128322 5918
rect 135438 5906 135490 5918
rect 122322 5854 122334 5906
rect 122386 5854 122398 5906
rect 124114 5854 124126 5906
rect 124178 5854 124190 5906
rect 129266 5854 129278 5906
rect 129330 5854 129342 5906
rect 130274 5854 130286 5906
rect 130338 5854 130350 5906
rect 134866 5854 134878 5906
rect 134930 5854 134942 5906
rect 119870 5842 119922 5854
rect 128270 5842 128322 5854
rect 135438 5842 135490 5854
rect 137342 5906 137394 5918
rect 140130 5854 140142 5906
rect 140194 5854 140206 5906
rect 141026 5854 141038 5906
rect 141090 5854 141102 5906
rect 142706 5854 142718 5906
rect 142770 5854 142782 5906
rect 145506 5854 145518 5906
rect 145570 5854 145582 5906
rect 137342 5842 137394 5854
rect 7982 5794 8034 5806
rect 7982 5730 8034 5742
rect 9662 5794 9714 5806
rect 9662 5730 9714 5742
rect 11230 5794 11282 5806
rect 11230 5730 11282 5742
rect 11790 5794 11842 5806
rect 11790 5730 11842 5742
rect 12686 5794 12738 5806
rect 12686 5730 12738 5742
rect 19854 5794 19906 5806
rect 31614 5794 31666 5806
rect 28578 5742 28590 5794
rect 28642 5742 28654 5794
rect 29922 5742 29934 5794
rect 29986 5742 29998 5794
rect 19854 5730 19906 5742
rect 31614 5730 31666 5742
rect 32062 5794 32114 5806
rect 40014 5794 40066 5806
rect 35074 5742 35086 5794
rect 35138 5742 35150 5794
rect 35634 5742 35646 5794
rect 35698 5742 35710 5794
rect 32062 5730 32114 5742
rect 40014 5730 40066 5742
rect 45054 5794 45106 5806
rect 45054 5730 45106 5742
rect 57934 5794 57986 5806
rect 57934 5730 57986 5742
rect 58606 5794 58658 5806
rect 58606 5730 58658 5742
rect 59502 5794 59554 5806
rect 65438 5794 65490 5806
rect 63746 5742 63758 5794
rect 63810 5742 63822 5794
rect 59502 5730 59554 5742
rect 65438 5730 65490 5742
rect 70926 5794 70978 5806
rect 74734 5794 74786 5806
rect 77086 5794 77138 5806
rect 71810 5742 71822 5794
rect 71874 5742 71886 5794
rect 76178 5742 76190 5794
rect 76242 5742 76254 5794
rect 70926 5730 70978 5742
rect 74734 5730 74786 5742
rect 77086 5730 77138 5742
rect 82462 5794 82514 5806
rect 90974 5794 91026 5806
rect 85586 5742 85598 5794
rect 85650 5742 85662 5794
rect 82462 5730 82514 5742
rect 90974 5730 91026 5742
rect 91758 5794 91810 5806
rect 91758 5730 91810 5742
rect 93998 5794 94050 5806
rect 93998 5730 94050 5742
rect 95790 5794 95842 5806
rect 106318 5794 106370 5806
rect 105410 5742 105422 5794
rect 105474 5742 105486 5794
rect 95790 5730 95842 5742
rect 106318 5730 106370 5742
rect 107326 5794 107378 5806
rect 113598 5794 113650 5806
rect 109890 5742 109902 5794
rect 109954 5742 109966 5794
rect 112130 5742 112142 5794
rect 112194 5742 112206 5794
rect 107326 5730 107378 5742
rect 113598 5730 113650 5742
rect 116510 5794 116562 5806
rect 121438 5794 121490 5806
rect 121090 5742 121102 5794
rect 121154 5742 121166 5794
rect 116510 5730 116562 5742
rect 121438 5730 121490 5742
rect 121998 5794 122050 5806
rect 121998 5730 122050 5742
rect 122110 5794 122162 5806
rect 125582 5794 125634 5806
rect 124002 5742 124014 5794
rect 124066 5742 124078 5794
rect 122110 5730 122162 5742
rect 125582 5730 125634 5742
rect 126030 5794 126082 5806
rect 126030 5730 126082 5742
rect 126478 5794 126530 5806
rect 126478 5730 126530 5742
rect 126814 5794 126866 5806
rect 126814 5730 126866 5742
rect 137790 5794 137842 5806
rect 137790 5730 137842 5742
rect 138910 5794 138962 5806
rect 138910 5730 138962 5742
rect 143950 5794 144002 5806
rect 143950 5730 144002 5742
rect 146078 5794 146130 5806
rect 146078 5730 146130 5742
rect 147310 5794 147362 5806
rect 147310 5730 147362 5742
rect 147758 5794 147810 5806
rect 147758 5730 147810 5742
rect 148206 5794 148258 5806
rect 148206 5730 148258 5742
rect 148766 5794 148818 5806
rect 148766 5730 148818 5742
rect 149102 5794 149154 5806
rect 149102 5730 149154 5742
rect 149662 5794 149714 5806
rect 149662 5730 149714 5742
rect 149998 5794 150050 5806
rect 149998 5730 150050 5742
rect 17838 5682 17890 5694
rect 17838 5618 17890 5630
rect 18174 5682 18226 5694
rect 43374 5682 43426 5694
rect 28914 5630 28926 5682
rect 28978 5679 28990 5682
rect 29474 5679 29486 5682
rect 28978 5633 29486 5679
rect 28978 5630 28990 5633
rect 29474 5630 29486 5633
rect 29538 5630 29550 5682
rect 18174 5618 18226 5630
rect 43374 5618 43426 5630
rect 68910 5682 68962 5694
rect 68910 5618 68962 5630
rect 92542 5682 92594 5694
rect 96014 5682 96066 5694
rect 103070 5682 103122 5694
rect 93314 5630 93326 5682
rect 93378 5679 93390 5682
rect 93986 5679 93998 5682
rect 93378 5633 93998 5679
rect 93378 5630 93390 5633
rect 93986 5630 93998 5633
rect 94050 5630 94062 5682
rect 97346 5630 97358 5682
rect 97410 5630 97422 5682
rect 101490 5630 101502 5682
rect 101554 5630 101566 5682
rect 92542 5618 92594 5630
rect 96014 5618 96066 5630
rect 103070 5618 103122 5630
rect 117742 5682 117794 5694
rect 117742 5618 117794 5630
rect 118526 5682 118578 5694
rect 118526 5618 118578 5630
rect 118750 5682 118802 5694
rect 118750 5618 118802 5630
rect 118862 5682 118914 5694
rect 118862 5618 118914 5630
rect 119422 5682 119474 5694
rect 119422 5618 119474 5630
rect 119534 5682 119586 5694
rect 127934 5682 127986 5694
rect 126018 5630 126030 5682
rect 126082 5679 126094 5682
rect 126242 5679 126254 5682
rect 126082 5633 126254 5679
rect 126082 5630 126094 5633
rect 126242 5630 126254 5633
rect 126306 5630 126318 5682
rect 126466 5630 126478 5682
rect 126530 5679 126542 5682
rect 126690 5679 126702 5682
rect 126530 5633 126702 5679
rect 126530 5630 126542 5633
rect 126690 5630 126702 5633
rect 126754 5630 126766 5682
rect 127026 5630 127038 5682
rect 127090 5679 127102 5682
rect 127362 5679 127374 5682
rect 127090 5633 127374 5679
rect 127090 5630 127102 5633
rect 127362 5630 127374 5633
rect 127426 5630 127438 5682
rect 119534 5618 119586 5630
rect 127934 5618 127986 5630
rect 129950 5682 130002 5694
rect 129950 5618 130002 5630
rect 130286 5682 130338 5694
rect 130286 5618 130338 5630
rect 133982 5682 134034 5694
rect 133982 5618 134034 5630
rect 139806 5682 139858 5694
rect 148642 5630 148654 5682
rect 148706 5679 148718 5682
rect 149090 5679 149102 5682
rect 148706 5633 149102 5679
rect 148706 5630 148718 5633
rect 149090 5630 149102 5633
rect 149154 5630 149166 5682
rect 139806 5618 139858 5630
rect 1344 5514 178640 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 96638 5514
rect 96690 5462 96742 5514
rect 96794 5462 96846 5514
rect 96898 5462 127358 5514
rect 127410 5462 127462 5514
rect 127514 5462 127566 5514
rect 127618 5462 158078 5514
rect 158130 5462 158182 5514
rect 158234 5462 158286 5514
rect 158338 5462 178640 5514
rect 1344 5428 178640 5462
rect 14590 5346 14642 5358
rect 8978 5294 8990 5346
rect 9042 5294 9054 5346
rect 14590 5282 14642 5294
rect 45950 5346 46002 5358
rect 45950 5282 46002 5294
rect 46286 5346 46338 5358
rect 46286 5282 46338 5294
rect 62302 5346 62354 5358
rect 62302 5282 62354 5294
rect 62638 5346 62690 5358
rect 69806 5346 69858 5358
rect 68450 5294 68462 5346
rect 68514 5294 68526 5346
rect 62638 5282 62690 5294
rect 69806 5282 69858 5294
rect 71374 5346 71426 5358
rect 71374 5282 71426 5294
rect 79998 5346 80050 5358
rect 79998 5282 80050 5294
rect 80894 5346 80946 5358
rect 80894 5282 80946 5294
rect 95902 5346 95954 5358
rect 95902 5282 95954 5294
rect 96238 5346 96290 5358
rect 96238 5282 96290 5294
rect 102062 5346 102114 5358
rect 110238 5346 110290 5358
rect 106754 5294 106766 5346
rect 106818 5343 106830 5346
rect 106978 5343 106990 5346
rect 106818 5297 106990 5343
rect 106818 5294 106830 5297
rect 106978 5294 106990 5297
rect 107042 5294 107054 5346
rect 102062 5282 102114 5294
rect 110238 5282 110290 5294
rect 111134 5346 111186 5358
rect 111134 5282 111186 5294
rect 111470 5346 111522 5358
rect 111470 5282 111522 5294
rect 119646 5346 119698 5358
rect 119646 5282 119698 5294
rect 123006 5346 123058 5358
rect 123006 5282 123058 5294
rect 123454 5346 123506 5358
rect 123454 5282 123506 5294
rect 123902 5346 123954 5358
rect 123902 5282 123954 5294
rect 125582 5346 125634 5358
rect 125582 5282 125634 5294
rect 125806 5346 125858 5358
rect 125806 5282 125858 5294
rect 133086 5346 133138 5358
rect 133086 5282 133138 5294
rect 133198 5346 133250 5358
rect 133198 5282 133250 5294
rect 133422 5346 133474 5358
rect 133422 5282 133474 5294
rect 136670 5346 136722 5358
rect 136670 5282 136722 5294
rect 136782 5346 136834 5358
rect 136782 5282 136834 5294
rect 137006 5346 137058 5358
rect 137006 5282 137058 5294
rect 137230 5346 137282 5358
rect 137230 5282 137282 5294
rect 139134 5346 139186 5358
rect 142942 5346 142994 5358
rect 139682 5294 139694 5346
rect 139746 5343 139758 5346
rect 139746 5297 139855 5343
rect 139746 5294 139758 5297
rect 139134 5282 139186 5294
rect 8430 5234 8482 5246
rect 8430 5170 8482 5182
rect 13694 5234 13746 5246
rect 21870 5234 21922 5246
rect 30718 5234 30770 5246
rect 36878 5234 36930 5246
rect 70030 5234 70082 5246
rect 75630 5234 75682 5246
rect 18946 5182 18958 5234
rect 19010 5182 19022 5234
rect 19842 5182 19854 5234
rect 19906 5182 19918 5234
rect 24098 5182 24110 5234
rect 24162 5182 24174 5234
rect 27794 5182 27806 5234
rect 27858 5182 27870 5234
rect 31490 5182 31502 5234
rect 31554 5182 31566 5234
rect 33058 5182 33070 5234
rect 33122 5182 33134 5234
rect 40450 5182 40462 5234
rect 40514 5182 40526 5234
rect 42578 5182 42590 5234
rect 42642 5182 42654 5234
rect 47394 5182 47406 5234
rect 47458 5182 47470 5234
rect 49746 5182 49758 5234
rect 49810 5182 49822 5234
rect 51874 5182 51886 5234
rect 51938 5182 51950 5234
rect 54562 5182 54574 5234
rect 54626 5182 54638 5234
rect 56690 5182 56702 5234
rect 56754 5182 56766 5234
rect 58482 5182 58494 5234
rect 58546 5182 58558 5234
rect 60610 5182 60622 5234
rect 60674 5182 60686 5234
rect 68226 5182 68238 5234
rect 68290 5182 68302 5234
rect 75282 5182 75294 5234
rect 75346 5182 75358 5234
rect 13694 5170 13746 5182
rect 21870 5170 21922 5182
rect 30718 5170 30770 5182
rect 36878 5170 36930 5182
rect 70030 5170 70082 5182
rect 75630 5170 75682 5182
rect 78206 5234 78258 5246
rect 78206 5170 78258 5182
rect 78654 5234 78706 5246
rect 84254 5234 84306 5246
rect 81218 5182 81230 5234
rect 81282 5182 81294 5234
rect 78654 5170 78706 5182
rect 84254 5170 84306 5182
rect 87390 5234 87442 5246
rect 87390 5170 87442 5182
rect 87502 5234 87554 5246
rect 87502 5170 87554 5182
rect 87614 5234 87666 5246
rect 87614 5170 87666 5182
rect 88174 5234 88226 5246
rect 91310 5234 91362 5246
rect 88946 5182 88958 5234
rect 89010 5182 89022 5234
rect 88174 5170 88226 5182
rect 91310 5170 91362 5182
rect 91646 5234 91698 5246
rect 91646 5170 91698 5182
rect 97806 5234 97858 5246
rect 97806 5170 97858 5182
rect 98030 5234 98082 5246
rect 98030 5170 98082 5182
rect 99598 5234 99650 5246
rect 99598 5170 99650 5182
rect 99822 5234 99874 5246
rect 99822 5170 99874 5182
rect 100270 5234 100322 5246
rect 100270 5170 100322 5182
rect 101054 5234 101106 5246
rect 101054 5170 101106 5182
rect 102286 5234 102338 5246
rect 102286 5170 102338 5182
rect 106318 5234 106370 5246
rect 106318 5170 106370 5182
rect 106654 5234 106706 5246
rect 119870 5234 119922 5246
rect 107762 5182 107774 5234
rect 107826 5182 107838 5234
rect 112242 5182 112254 5234
rect 112306 5182 112318 5234
rect 113810 5182 113822 5234
rect 113874 5182 113886 5234
rect 106654 5170 106706 5182
rect 119870 5170 119922 5182
rect 119982 5234 120034 5246
rect 119982 5170 120034 5182
rect 121662 5234 121714 5246
rect 121662 5170 121714 5182
rect 121774 5234 121826 5246
rect 121774 5170 121826 5182
rect 121886 5234 121938 5246
rect 121886 5170 121938 5182
rect 126030 5234 126082 5246
rect 126030 5170 126082 5182
rect 131742 5234 131794 5246
rect 131742 5170 131794 5182
rect 137790 5234 137842 5246
rect 137790 5170 137842 5182
rect 8654 5122 8706 5134
rect 7634 5070 7646 5122
rect 7698 5070 7710 5122
rect 8654 5058 8706 5070
rect 12014 5122 12066 5134
rect 12014 5058 12066 5070
rect 14254 5122 14306 5134
rect 37886 5122 37938 5134
rect 16146 5070 16158 5122
rect 16210 5070 16222 5122
rect 16818 5070 16830 5122
rect 16882 5070 16894 5122
rect 20738 5070 20750 5122
rect 20802 5070 20814 5122
rect 23426 5070 23438 5122
rect 23490 5070 23502 5122
rect 26898 5070 26910 5122
rect 26962 5070 26974 5122
rect 28690 5070 28702 5122
rect 28754 5070 28766 5122
rect 32274 5070 32286 5122
rect 32338 5070 32350 5122
rect 35970 5070 35982 5122
rect 36034 5070 36046 5122
rect 14254 5058 14306 5070
rect 37886 5058 37938 5070
rect 38222 5122 38274 5134
rect 43934 5122 43986 5134
rect 43250 5070 43262 5122
rect 43314 5070 43326 5122
rect 38222 5058 38274 5070
rect 43934 5058 43986 5070
rect 45390 5122 45442 5134
rect 66782 5122 66834 5134
rect 70254 5122 70306 5134
rect 77646 5122 77698 5134
rect 83582 5122 83634 5134
rect 48066 5070 48078 5122
rect 48130 5070 48142 5122
rect 52546 5070 52558 5122
rect 52610 5070 52622 5122
rect 53778 5070 53790 5122
rect 53842 5070 53854 5122
rect 57698 5070 57710 5122
rect 57762 5070 57774 5122
rect 61842 5070 61854 5122
rect 61906 5070 61918 5122
rect 66322 5070 66334 5122
rect 66386 5070 66398 5122
rect 67666 5070 67678 5122
rect 67730 5070 67742 5122
rect 72258 5070 72270 5122
rect 72322 5070 72334 5122
rect 73602 5070 73614 5122
rect 73666 5070 73678 5122
rect 81890 5070 81902 5122
rect 81954 5070 81966 5122
rect 45390 5058 45442 5070
rect 66782 5058 66834 5070
rect 70254 5058 70306 5070
rect 77646 5058 77698 5070
rect 83582 5058 83634 5070
rect 84478 5122 84530 5134
rect 84478 5058 84530 5070
rect 85486 5122 85538 5134
rect 85486 5058 85538 5070
rect 86718 5122 86770 5134
rect 90638 5122 90690 5134
rect 87154 5070 87166 5122
rect 87218 5070 87230 5122
rect 89058 5070 89070 5122
rect 89122 5070 89134 5122
rect 86718 5058 86770 5070
rect 90638 5058 90690 5070
rect 97134 5122 97186 5134
rect 98926 5122 98978 5134
rect 102510 5122 102562 5134
rect 104190 5122 104242 5134
rect 105646 5122 105698 5134
rect 109454 5122 109506 5134
rect 120094 5122 120146 5134
rect 98578 5070 98590 5122
rect 98642 5070 98654 5122
rect 101602 5070 101614 5122
rect 101666 5070 101678 5122
rect 103730 5070 103742 5122
rect 103794 5070 103806 5122
rect 105298 5070 105310 5122
rect 105362 5070 105374 5122
rect 107650 5070 107662 5122
rect 107714 5070 107726 5122
rect 110226 5070 110238 5122
rect 110290 5070 110302 5122
rect 112578 5070 112590 5122
rect 112642 5070 112654 5122
rect 113922 5070 113934 5122
rect 113986 5070 113998 5122
rect 115266 5070 115278 5122
rect 115330 5070 115342 5122
rect 119186 5070 119198 5122
rect 119250 5070 119262 5122
rect 97134 5058 97186 5070
rect 98926 5058 98978 5070
rect 102510 5058 102562 5070
rect 104190 5058 104242 5070
rect 105646 5058 105698 5070
rect 109454 5058 109506 5070
rect 120094 5058 120146 5070
rect 121214 5122 121266 5134
rect 121214 5058 121266 5070
rect 123678 5122 123730 5134
rect 123678 5058 123730 5070
rect 124910 5122 124962 5134
rect 124910 5058 124962 5070
rect 125358 5122 125410 5134
rect 125358 5058 125410 5070
rect 127262 5122 127314 5134
rect 127262 5058 127314 5070
rect 127710 5122 127762 5134
rect 127710 5058 127762 5070
rect 127934 5122 127986 5134
rect 127934 5058 127986 5070
rect 128158 5122 128210 5134
rect 128158 5058 128210 5070
rect 128382 5122 128434 5134
rect 128382 5058 128434 5070
rect 128942 5122 128994 5134
rect 128942 5058 128994 5070
rect 130510 5122 130562 5134
rect 130510 5058 130562 5070
rect 130734 5122 130786 5134
rect 130734 5058 130786 5070
rect 133646 5122 133698 5134
rect 133646 5058 133698 5070
rect 135998 5122 136050 5134
rect 139809 5122 139855 5297
rect 142942 5282 142994 5294
rect 143950 5346 144002 5358
rect 143950 5282 144002 5294
rect 147646 5234 147698 5246
rect 147646 5170 147698 5182
rect 143054 5122 143106 5134
rect 139794 5070 139806 5122
rect 139858 5070 139870 5122
rect 135998 5058 136050 5070
rect 143054 5058 143106 5070
rect 143278 5122 143330 5134
rect 143278 5058 143330 5070
rect 144062 5122 144114 5134
rect 152462 5122 152514 5134
rect 149090 5070 149102 5122
rect 149154 5070 149166 5122
rect 144062 5058 144114 5070
rect 152462 5058 152514 5070
rect 159294 5122 159346 5134
rect 159294 5058 159346 5070
rect 161086 5122 161138 5134
rect 161086 5058 161138 5070
rect 7870 5010 7922 5022
rect 7870 4946 7922 4958
rect 9550 5010 9602 5022
rect 9550 4946 9602 4958
rect 9886 5010 9938 5022
rect 9886 4946 9938 4958
rect 11230 5010 11282 5022
rect 11230 4946 11282 4958
rect 11566 5010 11618 5022
rect 11566 4946 11618 4958
rect 12910 5010 12962 5022
rect 30270 5010 30322 5022
rect 37550 5010 37602 5022
rect 14802 4958 14814 5010
rect 14866 4958 14878 5010
rect 15138 4958 15150 5010
rect 15202 4958 15214 5010
rect 22642 4958 22654 5010
rect 22706 4958 22718 5010
rect 26226 4958 26238 5010
rect 26290 4958 26302 5010
rect 35186 4958 35198 5010
rect 35250 4958 35262 5010
rect 12910 4946 12962 4958
rect 30270 4946 30322 4958
rect 37550 4946 37602 4958
rect 37998 5010 38050 5022
rect 37998 4946 38050 4958
rect 38670 5010 38722 5022
rect 38670 4946 38722 4958
rect 39006 5010 39058 5022
rect 39006 4946 39058 4958
rect 39566 5010 39618 5022
rect 39566 4946 39618 4958
rect 44382 5010 44434 5022
rect 44382 4946 44434 4958
rect 44718 5010 44770 5022
rect 44718 4946 44770 4958
rect 48862 5010 48914 5022
rect 48862 4946 48914 4958
rect 49198 5010 49250 5022
rect 64094 5010 64146 5022
rect 61506 4958 61518 5010
rect 61570 4958 61582 5010
rect 49198 4946 49250 4958
rect 64094 4946 64146 4958
rect 64430 5010 64482 5022
rect 64430 4946 64482 4958
rect 64990 5010 65042 5022
rect 64990 4946 65042 4958
rect 65326 5010 65378 5022
rect 65326 4946 65378 4958
rect 66894 5010 66946 5022
rect 66894 4946 66946 4958
rect 69358 5010 69410 5022
rect 70814 5010 70866 5022
rect 69570 4958 69582 5010
rect 69634 4958 69646 5010
rect 69358 4946 69410 4958
rect 70814 4946 70866 4958
rect 71038 5010 71090 5022
rect 71038 4946 71090 4958
rect 71262 5010 71314 5022
rect 76190 5010 76242 5022
rect 72482 4958 72494 5010
rect 72546 4958 72558 5010
rect 73490 4958 73502 5010
rect 73554 4958 73566 5010
rect 71262 4946 71314 4958
rect 76190 4946 76242 4958
rect 77982 5010 78034 5022
rect 77982 4946 78034 4958
rect 79102 5010 79154 5022
rect 79102 4946 79154 4958
rect 79438 5010 79490 5022
rect 79438 4946 79490 4958
rect 80222 5010 80274 5022
rect 80222 4946 80274 4958
rect 81118 5010 81170 5022
rect 81118 4946 81170 4958
rect 83470 5010 83522 5022
rect 83470 4946 83522 4958
rect 83918 5010 83970 5022
rect 83918 4946 83970 4958
rect 86494 5010 86546 5022
rect 86494 4946 86546 4958
rect 89742 5010 89794 5022
rect 89742 4946 89794 4958
rect 90414 5010 90466 5022
rect 90414 4946 90466 4958
rect 90974 5010 91026 5022
rect 90974 4946 91026 4958
rect 91422 5010 91474 5022
rect 91422 4946 91474 4958
rect 92430 5010 92482 5022
rect 92430 4946 92482 4958
rect 93214 5010 93266 5022
rect 93214 4946 93266 4958
rect 94110 5010 94162 5022
rect 94110 4946 94162 4958
rect 95006 5010 95058 5022
rect 95006 4946 95058 4958
rect 96126 5010 96178 5022
rect 96126 4946 96178 4958
rect 96910 5010 96962 5022
rect 96910 4946 96962 4958
rect 97470 5010 97522 5022
rect 97470 4946 97522 4958
rect 98814 5010 98866 5022
rect 98814 4946 98866 4958
rect 99262 5010 99314 5022
rect 102398 5010 102450 5022
rect 105982 5010 106034 5022
rect 101826 4958 101838 5010
rect 101890 4958 101902 5010
rect 103058 4958 103070 5010
rect 103122 4958 103134 5010
rect 104738 4958 104750 5010
rect 104802 4958 104814 5010
rect 99262 4946 99314 4958
rect 102398 4946 102450 4958
rect 105982 4946 106034 4958
rect 108334 5010 108386 5022
rect 108334 4946 108386 4958
rect 110574 5010 110626 5022
rect 110574 4946 110626 4958
rect 113038 5010 113090 5022
rect 113038 4946 113090 4958
rect 114606 5010 114658 5022
rect 114606 4946 114658 4958
rect 117070 5010 117122 5022
rect 117070 4946 117122 4958
rect 117406 5010 117458 5022
rect 117406 4946 117458 4958
rect 118302 5010 118354 5022
rect 118302 4946 118354 4958
rect 118638 5010 118690 5022
rect 120766 5010 120818 5022
rect 119410 4958 119422 5010
rect 119474 4958 119486 5010
rect 118638 4946 118690 4958
rect 120766 4946 120818 4958
rect 121326 5010 121378 5022
rect 121326 4946 121378 4958
rect 124126 5010 124178 5022
rect 124126 4946 124178 4958
rect 129278 5010 129330 5022
rect 129278 4946 129330 4958
rect 130622 5010 130674 5022
rect 130622 4946 130674 4958
rect 131070 5010 131122 5022
rect 131070 4946 131122 4958
rect 131630 5010 131682 5022
rect 131630 4946 131682 4958
rect 133758 5010 133810 5022
rect 133758 4946 133810 4958
rect 134318 5010 134370 5022
rect 134318 4946 134370 4958
rect 134654 5010 134706 5022
rect 134654 4946 134706 4958
rect 135438 5010 135490 5022
rect 135438 4946 135490 4958
rect 135662 5010 135714 5022
rect 135662 4946 135714 4958
rect 137342 5010 137394 5022
rect 137342 4946 137394 4958
rect 137902 5010 137954 5022
rect 137902 4946 137954 4958
rect 138350 5010 138402 5022
rect 138350 4946 138402 4958
rect 138574 5010 138626 5022
rect 138574 4946 138626 4958
rect 139358 5010 139410 5022
rect 139358 4946 139410 4958
rect 140926 5010 140978 5022
rect 140926 4946 140978 4958
rect 141262 5010 141314 5022
rect 141262 4946 141314 4958
rect 141822 5010 141874 5022
rect 141822 4946 141874 4958
rect 142158 5010 142210 5022
rect 142158 4946 142210 4958
rect 143390 5010 143442 5022
rect 143390 4946 143442 4958
rect 144958 5010 145010 5022
rect 144958 4946 145010 4958
rect 145294 5010 145346 5022
rect 145294 4946 145346 4958
rect 146190 5010 146242 5022
rect 146190 4946 146242 4958
rect 146750 5010 146802 5022
rect 146750 4946 146802 4958
rect 147086 5010 147138 5022
rect 147086 4946 147138 4958
rect 147758 5010 147810 5022
rect 147758 4946 147810 4958
rect 148878 5010 148930 5022
rect 148878 4946 148930 4958
rect 7086 4898 7138 4910
rect 7086 4834 7138 4846
rect 10782 4898 10834 4910
rect 10782 4834 10834 4846
rect 12574 4898 12626 4910
rect 12574 4834 12626 4846
rect 29934 4898 29986 4910
rect 29934 4834 29986 4846
rect 39902 4898 39954 4910
rect 39902 4834 39954 4846
rect 46174 4898 46226 4910
rect 46174 4834 46226 4846
rect 57262 4898 57314 4910
rect 57262 4834 57314 4846
rect 63646 4898 63698 4910
rect 76526 4898 76578 4910
rect 69682 4846 69694 4898
rect 69746 4846 69758 4898
rect 63646 4834 63698 4846
rect 76526 4834 76578 4846
rect 77422 4898 77474 4910
rect 77422 4834 77474 4846
rect 77534 4898 77586 4910
rect 77534 4834 77586 4846
rect 78094 4898 78146 4910
rect 78094 4834 78146 4846
rect 80110 4898 80162 4910
rect 80110 4834 80162 4846
rect 82126 4898 82178 4910
rect 82126 4834 82178 4846
rect 82686 4898 82738 4910
rect 82686 4834 82738 4846
rect 83358 4898 83410 4910
rect 83358 4834 83410 4846
rect 84030 4898 84082 4910
rect 84030 4834 84082 4846
rect 85822 4898 85874 4910
rect 85822 4834 85874 4846
rect 86606 4898 86658 4910
rect 86606 4834 86658 4846
rect 90526 4898 90578 4910
rect 90526 4834 90578 4846
rect 92094 4898 92146 4910
rect 92094 4834 92146 4846
rect 93550 4898 93602 4910
rect 93550 4834 93602 4846
rect 94446 4898 94498 4910
rect 94446 4834 94498 4846
rect 95342 4898 95394 4910
rect 95342 4834 95394 4846
rect 97022 4898 97074 4910
rect 97022 4834 97074 4846
rect 97582 4898 97634 4910
rect 97582 4834 97634 4846
rect 99374 4898 99426 4910
rect 105534 4898 105586 4910
rect 103618 4846 103630 4898
rect 103682 4846 103694 4898
rect 99374 4834 99426 4846
rect 105534 4834 105586 4846
rect 106094 4898 106146 4910
rect 106094 4834 106146 4846
rect 109118 4898 109170 4910
rect 109118 4834 109170 4846
rect 111358 4898 111410 4910
rect 111358 4834 111410 4846
rect 115502 4898 115554 4910
rect 115502 4834 115554 4846
rect 115950 4898 116002 4910
rect 115950 4834 116002 4846
rect 120878 4898 120930 4910
rect 120878 4834 120930 4846
rect 122446 4898 122498 4910
rect 122446 4834 122498 4846
rect 126590 4898 126642 4910
rect 126590 4834 126642 4846
rect 129838 4898 129890 4910
rect 129838 4834 129890 4846
rect 131854 4898 131906 4910
rect 131854 4834 131906 4846
rect 135886 4898 135938 4910
rect 135886 4834 135938 4846
rect 138126 4898 138178 4910
rect 138126 4834 138178 4846
rect 139246 4898 139298 4910
rect 139246 4834 139298 4846
rect 140030 4898 140082 4910
rect 140030 4834 140082 4846
rect 144174 4898 144226 4910
rect 144174 4834 144226 4846
rect 145854 4898 145906 4910
rect 145854 4834 145906 4846
rect 147870 4898 147922 4910
rect 147870 4834 147922 4846
rect 150110 4898 150162 4910
rect 150110 4834 150162 4846
rect 150670 4898 150722 4910
rect 150670 4834 150722 4846
rect 151230 4898 151282 4910
rect 151230 4834 151282 4846
rect 151790 4898 151842 4910
rect 151790 4834 151842 4846
rect 155374 4898 155426 4910
rect 155374 4834 155426 4846
rect 156718 4898 156770 4910
rect 156718 4834 156770 4846
rect 158398 4898 158450 4910
rect 158398 4834 158450 4846
rect 161534 4898 161586 4910
rect 161534 4834 161586 4846
rect 167134 4898 167186 4910
rect 167134 4834 167186 4846
rect 168030 4898 168082 4910
rect 168030 4834 168082 4846
rect 168926 4898 168978 4910
rect 168926 4834 168978 4846
rect 169374 4898 169426 4910
rect 169374 4834 169426 4846
rect 1344 4730 178640 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 81278 4730
rect 81330 4678 81382 4730
rect 81434 4678 81486 4730
rect 81538 4678 111998 4730
rect 112050 4678 112102 4730
rect 112154 4678 112206 4730
rect 112258 4678 142718 4730
rect 142770 4678 142822 4730
rect 142874 4678 142926 4730
rect 142978 4678 173438 4730
rect 173490 4678 173542 4730
rect 173594 4678 173646 4730
rect 173698 4678 178640 4730
rect 1344 4644 178640 4678
rect 10446 4562 10498 4574
rect 10446 4498 10498 4510
rect 16046 4562 16098 4574
rect 16046 4498 16098 4510
rect 16606 4562 16658 4574
rect 16606 4498 16658 4510
rect 18734 4562 18786 4574
rect 18734 4498 18786 4510
rect 23102 4562 23154 4574
rect 23102 4498 23154 4510
rect 26014 4562 26066 4574
rect 26014 4498 26066 4510
rect 26686 4562 26738 4574
rect 26686 4498 26738 4510
rect 33518 4562 33570 4574
rect 33518 4498 33570 4510
rect 39454 4562 39506 4574
rect 39454 4498 39506 4510
rect 40574 4562 40626 4574
rect 57822 4562 57874 4574
rect 40786 4510 40798 4562
rect 40850 4510 40862 4562
rect 40574 4498 40626 4510
rect 57822 4498 57874 4510
rect 61854 4562 61906 4574
rect 61854 4498 61906 4510
rect 62638 4562 62690 4574
rect 62638 4498 62690 4510
rect 64318 4562 64370 4574
rect 68910 4562 68962 4574
rect 67778 4510 67790 4562
rect 67842 4510 67854 4562
rect 64318 4498 64370 4510
rect 68910 4498 68962 4510
rect 71374 4562 71426 4574
rect 71374 4498 71426 4510
rect 72158 4562 72210 4574
rect 72158 4498 72210 4510
rect 74174 4562 74226 4574
rect 74174 4498 74226 4510
rect 78542 4562 78594 4574
rect 78542 4498 78594 4510
rect 78654 4562 78706 4574
rect 78654 4498 78706 4510
rect 81566 4562 81618 4574
rect 81566 4498 81618 4510
rect 83694 4562 83746 4574
rect 83694 4498 83746 4510
rect 84478 4562 84530 4574
rect 84478 4498 84530 4510
rect 84590 4562 84642 4574
rect 84590 4498 84642 4510
rect 85150 4562 85202 4574
rect 85150 4498 85202 4510
rect 90078 4562 90130 4574
rect 90078 4498 90130 4510
rect 90190 4562 90242 4574
rect 96350 4562 96402 4574
rect 91074 4510 91086 4562
rect 91138 4510 91150 4562
rect 93314 4510 93326 4562
rect 93378 4510 93390 4562
rect 90190 4498 90242 4510
rect 96350 4498 96402 4510
rect 100158 4562 100210 4574
rect 100158 4498 100210 4510
rect 100270 4562 100322 4574
rect 100270 4498 100322 4510
rect 100382 4562 100434 4574
rect 100382 4498 100434 4510
rect 101054 4562 101106 4574
rect 101054 4498 101106 4510
rect 102062 4562 102114 4574
rect 102062 4498 102114 4510
rect 105310 4562 105362 4574
rect 105310 4498 105362 4510
rect 105422 4562 105474 4574
rect 105422 4498 105474 4510
rect 108334 4562 108386 4574
rect 108334 4498 108386 4510
rect 109230 4562 109282 4574
rect 109230 4498 109282 4510
rect 113262 4562 113314 4574
rect 113262 4498 113314 4510
rect 113374 4562 113426 4574
rect 113374 4498 113426 4510
rect 113934 4562 113986 4574
rect 113934 4498 113986 4510
rect 114942 4562 114994 4574
rect 114942 4498 114994 4510
rect 115726 4562 115778 4574
rect 115726 4498 115778 4510
rect 116846 4562 116898 4574
rect 116846 4498 116898 4510
rect 117406 4562 117458 4574
rect 117406 4498 117458 4510
rect 117518 4562 117570 4574
rect 117518 4498 117570 4510
rect 118078 4562 118130 4574
rect 121326 4562 121378 4574
rect 122782 4562 122834 4574
rect 119746 4510 119758 4562
rect 119810 4510 119822 4562
rect 122210 4510 122222 4562
rect 122274 4510 122286 4562
rect 118078 4498 118130 4510
rect 121326 4498 121378 4510
rect 122782 4498 122834 4510
rect 123454 4562 123506 4574
rect 123454 4498 123506 4510
rect 123678 4562 123730 4574
rect 123678 4498 123730 4510
rect 124574 4562 124626 4574
rect 124574 4498 124626 4510
rect 126366 4562 126418 4574
rect 126366 4498 126418 4510
rect 127934 4562 127986 4574
rect 127934 4498 127986 4510
rect 133758 4562 133810 4574
rect 133758 4498 133810 4510
rect 135326 4562 135378 4574
rect 135326 4498 135378 4510
rect 138238 4562 138290 4574
rect 138238 4498 138290 4510
rect 139694 4562 139746 4574
rect 141710 4562 141762 4574
rect 141362 4510 141374 4562
rect 141426 4510 141438 4562
rect 139694 4498 139746 4510
rect 11454 4450 11506 4462
rect 39342 4450 39394 4462
rect 12786 4398 12798 4450
rect 12850 4398 12862 4450
rect 20066 4398 20078 4450
rect 20130 4398 20142 4450
rect 27570 4398 27582 4450
rect 27634 4398 27646 4450
rect 29922 4398 29934 4450
rect 29986 4398 29998 4450
rect 37986 4398 37998 4450
rect 38050 4398 38062 4450
rect 11454 4386 11506 4398
rect 39342 4386 39394 4398
rect 40126 4450 40178 4462
rect 43262 4450 43314 4462
rect 62302 4450 62354 4462
rect 42354 4398 42366 4450
rect 42418 4398 42430 4450
rect 47618 4398 47630 4450
rect 47682 4398 47694 4450
rect 51986 4398 51998 4450
rect 52050 4398 52062 4450
rect 60498 4398 60510 4450
rect 60562 4398 60574 4450
rect 40126 4386 40178 4398
rect 43262 4386 43314 4398
rect 62302 4386 62354 4398
rect 63198 4450 63250 4462
rect 63198 4386 63250 4398
rect 63534 4450 63586 4462
rect 63534 4386 63586 4398
rect 64430 4450 64482 4462
rect 68350 4450 68402 4462
rect 67666 4398 67678 4450
rect 67730 4398 67742 4450
rect 64430 4386 64482 4398
rect 68350 4386 68402 4398
rect 71822 4450 71874 4462
rect 71822 4386 71874 4398
rect 74062 4450 74114 4462
rect 74062 4386 74114 4398
rect 75630 4450 75682 4462
rect 75630 4386 75682 4398
rect 78430 4450 78482 4462
rect 78430 4386 78482 4398
rect 82014 4450 82066 4462
rect 82014 4386 82066 4398
rect 82350 4450 82402 4462
rect 82350 4386 82402 4398
rect 85038 4450 85090 4462
rect 85038 4386 85090 4398
rect 86382 4450 86434 4462
rect 86382 4386 86434 4398
rect 86718 4450 86770 4462
rect 86718 4386 86770 4398
rect 89294 4450 89346 4462
rect 89294 4386 89346 4398
rect 90638 4450 90690 4462
rect 90638 4386 90690 4398
rect 92094 4450 92146 4462
rect 92094 4386 92146 4398
rect 97358 4450 97410 4462
rect 97358 4386 97410 4398
rect 97470 4450 97522 4462
rect 97470 4386 97522 4398
rect 99822 4450 99874 4462
rect 99822 4386 99874 4398
rect 102958 4450 103010 4462
rect 102958 4386 103010 4398
rect 103294 4450 103346 4462
rect 103294 4386 103346 4398
rect 104414 4450 104466 4462
rect 104414 4386 104466 4398
rect 108894 4450 108946 4462
rect 108894 4386 108946 4398
rect 112030 4450 112082 4462
rect 112030 4386 112082 4398
rect 112366 4450 112418 4462
rect 112366 4386 112418 4398
rect 113822 4450 113874 4462
rect 113822 4386 113874 4398
rect 116174 4450 116226 4462
rect 116174 4386 116226 4398
rect 117966 4450 118018 4462
rect 117966 4386 118018 4398
rect 119422 4450 119474 4462
rect 120318 4450 120370 4462
rect 119634 4398 119646 4450
rect 119698 4398 119710 4450
rect 119422 4386 119474 4398
rect 120318 4386 120370 4398
rect 121774 4450 121826 4462
rect 121774 4386 121826 4398
rect 125582 4450 125634 4462
rect 125582 4386 125634 4398
rect 125806 4450 125858 4462
rect 125806 4386 125858 4398
rect 127822 4450 127874 4462
rect 127822 4386 127874 4398
rect 129054 4450 129106 4462
rect 129054 4386 129106 4398
rect 129278 4450 129330 4462
rect 129278 4386 129330 4398
rect 130062 4450 130114 4462
rect 130062 4386 130114 4398
rect 130286 4450 130338 4462
rect 130286 4386 130338 4398
rect 130846 4450 130898 4462
rect 130846 4386 130898 4398
rect 131070 4450 131122 4462
rect 131070 4386 131122 4398
rect 131742 4450 131794 4462
rect 131742 4386 131794 4398
rect 131966 4450 132018 4462
rect 131966 4386 132018 4398
rect 132974 4450 133026 4462
rect 133870 4450 133922 4462
rect 133186 4398 133198 4450
rect 133250 4447 133262 4450
rect 133410 4447 133422 4450
rect 133250 4401 133422 4447
rect 133250 4398 133262 4401
rect 133410 4398 133422 4401
rect 133474 4398 133486 4450
rect 132974 4386 133026 4398
rect 133870 4386 133922 4398
rect 134766 4450 134818 4462
rect 134766 4386 134818 4398
rect 135662 4450 135714 4462
rect 135662 4386 135714 4398
rect 136110 4450 136162 4462
rect 136110 4386 136162 4398
rect 137006 4450 137058 4462
rect 137006 4386 137058 4398
rect 139582 4450 139634 4462
rect 139582 4386 139634 4398
rect 139806 4450 139858 4462
rect 139806 4386 139858 4398
rect 140366 4450 140418 4462
rect 140366 4386 140418 4398
rect 10110 4338 10162 4350
rect 16942 4338 16994 4350
rect 8530 4286 8542 4338
rect 8594 4286 8606 4338
rect 11218 4286 11230 4338
rect 11282 4286 11294 4338
rect 12114 4286 12126 4338
rect 12178 4286 12190 4338
rect 15810 4286 15822 4338
rect 15874 4286 15886 4338
rect 10110 4274 10162 4286
rect 16942 4274 16994 4286
rect 18398 4338 18450 4350
rect 27022 4338 27074 4350
rect 32846 4338 32898 4350
rect 39678 4338 39730 4350
rect 19282 4286 19294 4338
rect 19346 4286 19358 4338
rect 22866 4286 22878 4338
rect 22930 4286 22942 4338
rect 23762 4286 23774 4338
rect 23826 4286 23838 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 27458 4286 27470 4338
rect 27522 4286 27534 4338
rect 29138 4286 29150 4338
rect 29202 4286 29214 4338
rect 34290 4286 34302 4338
rect 34354 4286 34366 4338
rect 38658 4286 38670 4338
rect 38722 4286 38734 4338
rect 18398 4274 18450 4286
rect 27022 4274 27074 4286
rect 32846 4274 32898 4286
rect 39678 4274 39730 4286
rect 40350 4338 40402 4350
rect 40350 4274 40402 4286
rect 40798 4338 40850 4350
rect 40798 4274 40850 4286
rect 42254 4338 42306 4350
rect 42254 4274 42306 4286
rect 42590 4338 42642 4350
rect 57486 4338 57538 4350
rect 67342 4338 67394 4350
rect 42802 4286 42814 4338
rect 42866 4286 42878 4338
rect 44930 4286 44942 4338
rect 44994 4286 45006 4338
rect 48402 4286 48414 4338
rect 48466 4286 48478 4338
rect 53890 4286 53902 4338
rect 53954 4286 53966 4338
rect 56578 4286 56590 4338
rect 56642 4286 56654 4338
rect 61170 4286 61182 4338
rect 61234 4286 61246 4338
rect 64082 4286 64094 4338
rect 64146 4286 64158 4338
rect 65538 4286 65550 4338
rect 65602 4286 65614 4338
rect 42590 4274 42642 4286
rect 57486 4274 57538 4286
rect 67342 4274 67394 4286
rect 67902 4338 67954 4350
rect 67902 4274 67954 4286
rect 68126 4338 68178 4350
rect 71710 4338 71762 4350
rect 69346 4286 69358 4338
rect 69410 4286 69422 4338
rect 71138 4286 71150 4338
rect 71202 4286 71214 4338
rect 68126 4274 68178 4286
rect 71710 4274 71762 4286
rect 72382 4338 72434 4350
rect 73614 4338 73666 4350
rect 73378 4286 73390 4338
rect 73442 4286 73454 4338
rect 72382 4274 72434 4286
rect 73614 4274 73666 4286
rect 73726 4338 73778 4350
rect 73726 4274 73778 4286
rect 74398 4338 74450 4350
rect 82798 4338 82850 4350
rect 75394 4286 75406 4338
rect 75458 4286 75470 4338
rect 76178 4286 76190 4338
rect 76242 4286 76254 4338
rect 79314 4286 79326 4338
rect 79378 4286 79390 4338
rect 74398 4274 74450 4286
rect 82798 4274 82850 4286
rect 83246 4338 83298 4350
rect 83246 4274 83298 4286
rect 83358 4338 83410 4350
rect 83358 4274 83410 4286
rect 83582 4338 83634 4350
rect 83582 4274 83634 4286
rect 83806 4338 83858 4350
rect 83806 4274 83858 4286
rect 84702 4338 84754 4350
rect 84702 4274 84754 4286
rect 85374 4338 85426 4350
rect 85374 4274 85426 4286
rect 85598 4338 85650 4350
rect 89406 4338 89458 4350
rect 88274 4286 88286 4338
rect 88338 4286 88350 4338
rect 85598 4274 85650 4286
rect 89406 4274 89458 4286
rect 90302 4338 90354 4350
rect 90302 4274 90354 4286
rect 91198 4338 91250 4350
rect 91198 4274 91250 4286
rect 91758 4338 91810 4350
rect 91758 4274 91810 4286
rect 92766 4338 92818 4350
rect 92766 4274 92818 4286
rect 92990 4338 93042 4350
rect 100046 4338 100098 4350
rect 94658 4286 94670 4338
rect 94722 4286 94734 4338
rect 98242 4286 98254 4338
rect 98306 4286 98318 4338
rect 92990 4274 93042 4286
rect 100046 4274 100098 4286
rect 101166 4338 101218 4350
rect 101950 4338 102002 4350
rect 101714 4286 101726 4338
rect 101778 4286 101790 4338
rect 101166 4274 101218 4286
rect 101950 4274 102002 4286
rect 102174 4338 102226 4350
rect 105982 4338 106034 4350
rect 108446 4338 108498 4350
rect 102386 4286 102398 4338
rect 102450 4286 102462 4338
rect 104178 4286 104190 4338
rect 104242 4286 104254 4338
rect 105634 4286 105646 4338
rect 105698 4286 105710 4338
rect 106530 4286 106542 4338
rect 106594 4286 106606 4338
rect 102174 4274 102226 4286
rect 105982 4274 106034 4286
rect 108446 4274 108498 4286
rect 108558 4338 108610 4350
rect 108558 4274 108610 4286
rect 109230 4338 109282 4350
rect 113710 4338 113762 4350
rect 111010 4286 111022 4338
rect 111074 4286 111086 4338
rect 109230 4274 109282 4286
rect 113710 4274 113762 4286
rect 114158 4338 114210 4350
rect 116062 4338 116114 4350
rect 115490 4286 115502 4338
rect 115554 4286 115566 4338
rect 114158 4274 114210 4286
rect 116062 4274 116114 4286
rect 116510 4338 116562 4350
rect 116510 4274 116562 4286
rect 116734 4338 116786 4350
rect 116734 4274 116786 4286
rect 117630 4338 117682 4350
rect 117630 4274 117682 4286
rect 119870 4338 119922 4350
rect 119870 4274 119922 4286
rect 121214 4338 121266 4350
rect 121214 4274 121266 4286
rect 121438 4338 121490 4350
rect 121438 4274 121490 4286
rect 122110 4338 122162 4350
rect 122110 4274 122162 4286
rect 122334 4338 122386 4350
rect 126702 4338 126754 4350
rect 124002 4286 124014 4338
rect 124066 4286 124078 4338
rect 124786 4286 124798 4338
rect 124850 4286 124862 4338
rect 122334 4274 122386 4286
rect 126702 4274 126754 4286
rect 132638 4338 132690 4350
rect 137342 4338 137394 4350
rect 138350 4338 138402 4350
rect 133522 4286 133534 4338
rect 133586 4286 133598 4338
rect 134418 4286 134430 4338
rect 134482 4286 134494 4338
rect 137554 4286 137566 4338
rect 137618 4286 137630 4338
rect 138114 4286 138126 4338
rect 138178 4286 138190 4338
rect 132638 4274 132690 4286
rect 137342 4274 137394 4286
rect 138350 4274 138402 4286
rect 138798 4338 138850 4350
rect 140578 4286 140590 4338
rect 140642 4286 140654 4338
rect 138798 4274 138850 4286
rect 6862 4226 6914 4238
rect 9102 4226 9154 4238
rect 17838 4226 17890 4238
rect 28590 4226 28642 4238
rect 41694 4226 41746 4238
rect 72046 4226 72098 4238
rect 7522 4174 7534 4226
rect 7586 4174 7598 4226
rect 14914 4174 14926 4226
rect 14978 4174 14990 4226
rect 22194 4174 22206 4226
rect 22258 4174 22270 4226
rect 24434 4174 24446 4226
rect 24498 4174 24510 4226
rect 32050 4174 32062 4226
rect 32114 4174 32126 4226
rect 34738 4174 34750 4226
rect 34802 4174 34814 4226
rect 35858 4174 35870 4226
rect 35922 4174 35934 4226
rect 44258 4174 44270 4226
rect 44322 4174 44334 4226
rect 45490 4174 45502 4226
rect 45554 4174 45566 4226
rect 55570 4174 55582 4226
rect 55634 4174 55646 4226
rect 58370 4174 58382 4226
rect 58434 4174 58446 4226
rect 66098 4174 66110 4226
rect 66162 4174 66174 4226
rect 70018 4174 70030 4226
rect 70082 4174 70094 4226
rect 6862 4162 6914 4174
rect 9102 4162 9154 4174
rect 17838 4162 17890 4174
rect 28590 4162 28642 4174
rect 41694 4162 41746 4174
rect 72046 4162 72098 4174
rect 74622 4226 74674 4238
rect 77982 4226 78034 4238
rect 90974 4226 91026 4238
rect 76850 4174 76862 4226
rect 76914 4174 76926 4226
rect 79986 4174 79998 4226
rect 80050 4174 80062 4226
rect 87714 4174 87726 4226
rect 87778 4174 87790 4226
rect 74622 4162 74674 4174
rect 77982 4162 78034 4174
rect 90974 4162 91026 4174
rect 93774 4226 93826 4238
rect 109454 4226 109506 4238
rect 114494 4226 114546 4238
rect 95330 4174 95342 4226
rect 95394 4174 95406 4226
rect 98690 4174 98702 4226
rect 98754 4174 98766 4226
rect 107090 4174 107102 4226
rect 107154 4174 107166 4226
rect 110226 4174 110238 4226
rect 110290 4174 110302 4226
rect 93774 4162 93826 4174
rect 109454 4162 109506 4174
rect 114494 4162 114546 4174
rect 118190 4226 118242 4238
rect 118190 4162 118242 4174
rect 118638 4226 118690 4238
rect 118638 4162 118690 4174
rect 120094 4226 120146 4238
rect 120094 4162 120146 4174
rect 123566 4226 123618 4238
rect 127150 4226 127202 4238
rect 125458 4174 125470 4226
rect 125522 4174 125534 4226
rect 123566 4162 123618 4174
rect 127150 4162 127202 4174
rect 129166 4226 129218 4238
rect 137118 4226 137170 4238
rect 129938 4174 129950 4226
rect 130002 4174 130014 4226
rect 131170 4174 131182 4226
rect 131234 4174 131246 4226
rect 132066 4174 132078 4226
rect 132130 4174 132142 4226
rect 134530 4174 134542 4226
rect 134594 4174 134606 4226
rect 129166 4162 129218 4174
rect 137118 4162 137170 4174
rect 128046 4114 128098 4126
rect 128046 4050 128098 4062
rect 138574 4114 138626 4126
rect 141377 4114 141423 4510
rect 141710 4498 141762 4510
rect 144062 4562 144114 4574
rect 144062 4498 144114 4510
rect 146078 4562 146130 4574
rect 146078 4498 146130 4510
rect 151230 4562 151282 4574
rect 151230 4498 151282 4510
rect 156270 4562 156322 4574
rect 156270 4498 156322 4510
rect 159070 4562 159122 4574
rect 159070 4498 159122 4510
rect 161310 4562 161362 4574
rect 161310 4498 161362 4510
rect 144958 4450 145010 4462
rect 144958 4386 145010 4398
rect 145518 4450 145570 4462
rect 145518 4386 145570 4398
rect 146974 4450 147026 4462
rect 146974 4386 147026 4398
rect 147870 4450 147922 4462
rect 147870 4386 147922 4398
rect 148094 4450 148146 4462
rect 148094 4386 148146 4398
rect 149662 4450 149714 4462
rect 149662 4386 149714 4398
rect 149998 4450 150050 4462
rect 149998 4386 150050 4398
rect 150558 4450 150610 4462
rect 150558 4386 150610 4398
rect 153470 4450 153522 4462
rect 153470 4386 153522 4398
rect 155150 4450 155202 4462
rect 155150 4386 155202 4398
rect 157166 4450 157218 4462
rect 157166 4386 157218 4398
rect 158398 4450 158450 4462
rect 158398 4386 158450 4398
rect 159966 4450 160018 4462
rect 159966 4386 160018 4398
rect 162206 4450 162258 4462
rect 162206 4386 162258 4398
rect 163550 4450 163602 4462
rect 163550 4386 163602 4398
rect 165230 4450 165282 4462
rect 165230 4386 165282 4398
rect 166910 4450 166962 4462
rect 166910 4386 166962 4398
rect 168030 4450 168082 4462
rect 168030 4386 168082 4398
rect 169150 4450 169202 4462
rect 169150 4386 169202 4398
rect 170270 4450 170322 4462
rect 170270 4386 170322 4398
rect 171950 4450 172002 4462
rect 171950 4386 172002 4398
rect 173070 4450 173122 4462
rect 173070 4386 173122 4398
rect 141822 4338 141874 4350
rect 141586 4286 141598 4338
rect 141650 4286 141662 4338
rect 141822 4274 141874 4286
rect 142046 4338 142098 4350
rect 142046 4274 142098 4286
rect 142830 4338 142882 4350
rect 142830 4274 142882 4286
rect 143278 4338 143330 4350
rect 143278 4274 143330 4286
rect 143502 4338 143554 4350
rect 143502 4274 143554 4286
rect 145070 4338 145122 4350
rect 145070 4274 145122 4286
rect 145182 4338 145234 4350
rect 148766 4338 148818 4350
rect 146290 4286 146302 4338
rect 146354 4286 146366 4338
rect 147298 4286 147310 4338
rect 147362 4286 147374 4338
rect 149090 4286 149102 4338
rect 149154 4286 149166 4338
rect 151442 4286 151454 4338
rect 151506 4286 151518 4338
rect 156482 4286 156494 4338
rect 156546 4286 156558 4338
rect 161522 4286 161534 4338
rect 161586 4286 161598 4338
rect 169362 4286 169374 4338
rect 169426 4286 169438 4338
rect 145182 4274 145234 4286
rect 148766 4274 148818 4286
rect 142270 4226 142322 4238
rect 142270 4162 142322 4174
rect 143054 4226 143106 4238
rect 143054 4162 143106 4174
rect 144174 4226 144226 4238
rect 152014 4226 152066 4238
rect 148978 4174 148990 4226
rect 149042 4174 149054 4226
rect 144174 4162 144226 4174
rect 152014 4162 152066 4174
rect 152798 4226 152850 4238
rect 152798 4162 152850 4174
rect 154030 4226 154082 4238
rect 154030 4162 154082 4174
rect 154590 4226 154642 4238
rect 154590 4162 154642 4174
rect 155822 4226 155874 4238
rect 155822 4162 155874 4174
rect 157726 4226 157778 4238
rect 157726 4162 157778 4174
rect 159182 4226 159234 4238
rect 159182 4162 159234 4174
rect 160750 4226 160802 4238
rect 160750 4162 160802 4174
rect 162766 4226 162818 4238
rect 162766 4162 162818 4174
rect 164110 4226 164162 4238
rect 164110 4162 164162 4174
rect 164558 4226 164610 4238
rect 164558 4162 164610 4174
rect 165790 4226 165842 4238
rect 165790 4162 165842 4174
rect 166350 4226 166402 4238
rect 166350 4162 166402 4174
rect 170830 4226 170882 4238
rect 170830 4162 170882 4174
rect 171390 4226 171442 4238
rect 171390 4162 171442 4174
rect 172510 4226 172562 4238
rect 172510 4162 172562 4174
rect 173630 4226 173682 4238
rect 173630 4162 173682 4174
rect 147310 4114 147362 4126
rect 141362 4062 141374 4114
rect 141426 4062 141438 4114
rect 138574 4050 138626 4062
rect 147310 4050 147362 4062
rect 148206 4114 148258 4126
rect 148206 4050 148258 4062
rect 1344 3946 178640 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 96638 3946
rect 96690 3894 96742 3946
rect 96794 3894 96846 3946
rect 96898 3894 127358 3946
rect 127410 3894 127462 3946
rect 127514 3894 127566 3946
rect 127618 3894 158078 3946
rect 158130 3894 158182 3946
rect 158234 3894 158286 3946
rect 158338 3894 178640 3946
rect 1344 3860 178640 3894
rect 21534 3778 21586 3790
rect 21534 3714 21586 3726
rect 21870 3778 21922 3790
rect 21870 3714 21922 3726
rect 26350 3778 26402 3790
rect 26350 3714 26402 3726
rect 26686 3778 26738 3790
rect 26686 3714 26738 3726
rect 30382 3778 30434 3790
rect 30382 3714 30434 3726
rect 30718 3778 30770 3790
rect 76974 3778 77026 3790
rect 64306 3726 64318 3778
rect 64370 3775 64382 3778
rect 64978 3775 64990 3778
rect 64370 3729 64990 3775
rect 64370 3726 64382 3729
rect 64978 3726 64990 3729
rect 65042 3726 65054 3778
rect 30718 3714 30770 3726
rect 76974 3714 77026 3726
rect 13806 3666 13858 3678
rect 8306 3614 8318 3666
rect 8370 3614 8382 3666
rect 10322 3614 10334 3666
rect 10386 3614 10398 3666
rect 12562 3614 12574 3666
rect 12626 3614 12638 3666
rect 13806 3602 13858 3614
rect 32510 3666 32562 3678
rect 64766 3666 64818 3678
rect 76526 3666 76578 3678
rect 37874 3614 37886 3666
rect 37938 3614 37950 3666
rect 39554 3614 39566 3666
rect 39618 3614 39630 3666
rect 41794 3614 41806 3666
rect 41858 3614 41870 3666
rect 43138 3614 43150 3666
rect 43202 3614 43214 3666
rect 49074 3614 49086 3666
rect 49138 3614 49150 3666
rect 51202 3614 51214 3666
rect 51266 3614 51278 3666
rect 53106 3614 53118 3666
rect 53170 3614 53182 3666
rect 61394 3614 61406 3666
rect 61458 3614 61470 3666
rect 63074 3614 63086 3666
rect 63138 3614 63150 3666
rect 71026 3614 71038 3666
rect 71090 3614 71102 3666
rect 72706 3614 72718 3666
rect 72770 3614 72782 3666
rect 32510 3602 32562 3614
rect 64766 3602 64818 3614
rect 76526 3602 76578 3614
rect 77086 3666 77138 3678
rect 88286 3666 88338 3678
rect 80994 3614 81006 3666
rect 81058 3614 81070 3666
rect 82786 3614 82798 3666
rect 82850 3614 82862 3666
rect 86258 3614 86270 3666
rect 86322 3614 86334 3666
rect 77086 3602 77138 3614
rect 88286 3602 88338 3614
rect 88734 3666 88786 3678
rect 88734 3602 88786 3614
rect 89182 3666 89234 3678
rect 89182 3602 89234 3614
rect 95790 3666 95842 3678
rect 95790 3602 95842 3614
rect 98926 3666 98978 3678
rect 109902 3666 109954 3678
rect 104962 3614 104974 3666
rect 105026 3663 105038 3666
rect 105522 3663 105534 3666
rect 105026 3617 105534 3663
rect 105026 3614 105038 3617
rect 105522 3614 105534 3617
rect 105586 3614 105598 3666
rect 98926 3602 98978 3614
rect 109902 3602 109954 3614
rect 110350 3666 110402 3678
rect 129950 3666 130002 3678
rect 114034 3614 114046 3666
rect 114098 3614 114110 3666
rect 117954 3614 117966 3666
rect 118018 3614 118030 3666
rect 121762 3614 121774 3666
rect 121826 3614 121838 3666
rect 110350 3602 110402 3614
rect 129950 3602 130002 3614
rect 148766 3666 148818 3678
rect 148766 3602 148818 3614
rect 14254 3554 14306 3566
rect 65214 3554 65266 3566
rect 98478 3554 98530 3566
rect 107550 3554 107602 3566
rect 110798 3554 110850 3566
rect 121438 3554 121490 3566
rect 6514 3502 6526 3554
rect 6578 3502 6590 3554
rect 10770 3502 10782 3554
rect 10834 3502 10846 3554
rect 11666 3502 11678 3554
rect 11730 3502 11742 3554
rect 15138 3502 15150 3554
rect 15202 3502 15214 3554
rect 18722 3502 18734 3554
rect 18786 3502 18798 3554
rect 20626 3502 20638 3554
rect 20690 3502 20702 3554
rect 22530 3502 22542 3554
rect 22594 3502 22606 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 25442 3502 25454 3554
rect 25506 3502 25518 3554
rect 27458 3502 27470 3554
rect 27522 3502 27534 3554
rect 28242 3502 28254 3554
rect 28306 3502 28318 3554
rect 29474 3502 29486 3554
rect 29538 3502 29550 3554
rect 34402 3502 34414 3554
rect 34466 3502 34478 3554
rect 36306 3502 36318 3554
rect 36370 3502 36382 3554
rect 37426 3502 37438 3554
rect 37490 3502 37502 3554
rect 40226 3502 40238 3554
rect 40290 3502 40302 3554
rect 41122 3502 41134 3554
rect 41186 3502 41198 3554
rect 44034 3502 44046 3554
rect 44098 3502 44110 3554
rect 46050 3502 46062 3554
rect 46114 3502 46126 3554
rect 46834 3502 46846 3554
rect 46898 3502 46910 3554
rect 51986 3502 51998 3554
rect 52050 3502 52062 3554
rect 54114 3502 54126 3554
rect 54178 3502 54190 3554
rect 55682 3502 55694 3554
rect 55746 3502 55758 3554
rect 57922 3502 57934 3554
rect 57986 3502 57998 3554
rect 59826 3502 59838 3554
rect 59890 3502 59902 3554
rect 60834 3502 60846 3554
rect 60898 3502 60910 3554
rect 63522 3502 63534 3554
rect 63586 3502 63598 3554
rect 66098 3502 66110 3554
rect 66162 3502 66174 3554
rect 68450 3502 68462 3554
rect 68514 3502 68526 3554
rect 70354 3502 70366 3554
rect 70418 3502 70430 3554
rect 73714 3502 73726 3554
rect 73778 3502 73790 3554
rect 74274 3502 74286 3554
rect 74338 3502 74350 3554
rect 77298 3502 77310 3554
rect 77362 3502 77374 3554
rect 77858 3502 77870 3554
rect 77922 3502 77934 3554
rect 80322 3502 80334 3554
rect 80386 3502 80398 3554
rect 82114 3502 82126 3554
rect 82178 3502 82190 3554
rect 84242 3502 84254 3554
rect 84306 3502 84318 3554
rect 87042 3502 87054 3554
rect 87106 3502 87118 3554
rect 89618 3502 89630 3554
rect 89682 3502 89694 3554
rect 92082 3502 92094 3554
rect 92146 3502 92158 3554
rect 93762 3502 93774 3554
rect 93826 3502 93838 3554
rect 94658 3502 94670 3554
rect 94722 3502 94734 3554
rect 96450 3502 96462 3554
rect 96514 3502 96526 3554
rect 99922 3502 99934 3554
rect 99986 3502 99998 3554
rect 102834 3502 102846 3554
rect 102898 3502 102910 3554
rect 104738 3502 104750 3554
rect 104802 3502 104814 3554
rect 105522 3502 105534 3554
rect 105586 3502 105598 3554
rect 108210 3502 108222 3554
rect 108274 3502 108286 3554
rect 112802 3502 112814 3554
rect 112866 3502 112878 3554
rect 113362 3502 113374 3554
rect 113426 3502 113438 3554
rect 115714 3502 115726 3554
rect 115778 3502 115790 3554
rect 117282 3502 117294 3554
rect 117346 3502 117358 3554
rect 119410 3502 119422 3554
rect 119474 3502 119486 3554
rect 121202 3502 121214 3554
rect 121266 3502 121278 3554
rect 14254 3490 14306 3502
rect 65214 3490 65266 3502
rect 98478 3490 98530 3502
rect 107550 3490 107602 3502
rect 110798 3490 110850 3502
rect 121438 3490 121490 3502
rect 121662 3554 121714 3566
rect 121662 3490 121714 3502
rect 123678 3554 123730 3566
rect 126366 3554 126418 3566
rect 124450 3502 124462 3554
rect 124514 3502 124526 3554
rect 125346 3502 125358 3554
rect 125410 3502 125422 3554
rect 123678 3490 123730 3502
rect 126366 3490 126418 3502
rect 127262 3554 127314 3566
rect 127262 3490 127314 3502
rect 128494 3554 128546 3566
rect 128494 3490 128546 3502
rect 129054 3554 129106 3566
rect 129054 3490 129106 3502
rect 131518 3554 131570 3566
rect 131518 3490 131570 3502
rect 132078 3554 132130 3566
rect 132078 3490 132130 3502
rect 134206 3554 134258 3566
rect 134206 3490 134258 3502
rect 135438 3554 135490 3566
rect 139022 3554 139074 3566
rect 137106 3502 137118 3554
rect 137170 3502 137182 3554
rect 138002 3502 138014 3554
rect 138066 3502 138078 3554
rect 135438 3490 135490 3502
rect 139022 3490 139074 3502
rect 140254 3554 140306 3566
rect 140254 3490 140306 3502
rect 141150 3554 141202 3566
rect 141150 3490 141202 3502
rect 143278 3554 143330 3566
rect 143278 3490 143330 3502
rect 144174 3554 144226 3566
rect 147198 3554 147250 3566
rect 144946 3502 144958 3554
rect 145010 3502 145022 3554
rect 144174 3490 144226 3502
rect 147198 3490 147250 3502
rect 148094 3554 148146 3566
rect 149886 3554 149938 3566
rect 148978 3502 148990 3554
rect 149042 3502 149054 3554
rect 148094 3490 148146 3502
rect 149886 3490 149938 3502
rect 151118 3554 151170 3566
rect 158958 3554 159010 3566
rect 161646 3554 161698 3566
rect 169486 3554 169538 3566
rect 151890 3502 151902 3554
rect 151954 3502 151966 3554
rect 153682 3502 153694 3554
rect 153746 3502 153758 3554
rect 155810 3502 155822 3554
rect 155874 3502 155886 3554
rect 156706 3502 156718 3554
rect 156770 3502 156782 3554
rect 157602 3502 157614 3554
rect 157666 3502 157678 3554
rect 160626 3502 160638 3554
rect 160690 3502 160702 3554
rect 163650 3502 163662 3554
rect 163714 3502 163726 3554
rect 165442 3502 165454 3554
rect 165506 3502 165518 3554
rect 167570 3502 167582 3554
rect 167634 3502 167646 3554
rect 151118 3490 151170 3502
rect 158958 3490 159010 3502
rect 161646 3490 161698 3502
rect 169486 3490 169538 3502
rect 170718 3554 170770 3566
rect 173406 3554 173458 3566
rect 172386 3502 172398 3554
rect 172450 3502 172462 3554
rect 170718 3490 170770 3502
rect 173406 3490 173458 3502
rect 5854 3442 5906 3454
rect 121774 3442 121826 3454
rect 16034 3390 16046 3442
rect 16098 3390 16110 3442
rect 17826 3390 17838 3442
rect 17890 3390 17902 3442
rect 19730 3390 19742 3442
rect 19794 3390 19806 3442
rect 22418 3390 22430 3442
rect 22482 3390 22494 3442
rect 23650 3390 23662 3442
rect 23714 3390 23726 3442
rect 27234 3390 27246 3442
rect 27298 3390 27310 3442
rect 30930 3390 30942 3442
rect 30994 3390 31006 3442
rect 31490 3390 31502 3442
rect 31554 3390 31566 3442
rect 33506 3390 33518 3442
rect 33570 3390 33582 3442
rect 35410 3390 35422 3442
rect 35474 3390 35486 3442
rect 45378 3390 45390 3442
rect 45442 3390 45454 3442
rect 47730 3390 47742 3442
rect 47794 3390 47806 3442
rect 55010 3390 55022 3442
rect 55074 3390 55086 3442
rect 57138 3390 57150 3442
rect 57202 3390 57214 3442
rect 58930 3390 58942 3442
rect 58994 3390 59006 3442
rect 66994 3390 67006 3442
rect 67058 3390 67070 3442
rect 69346 3390 69358 3442
rect 69410 3390 69422 3442
rect 75170 3390 75182 3442
rect 75234 3390 75246 3442
rect 78754 3390 78766 3442
rect 78818 3390 78830 3442
rect 85138 3390 85150 3442
rect 85202 3390 85214 3442
rect 90514 3390 90526 3442
rect 90578 3390 90590 3442
rect 92866 3390 92878 3442
rect 92930 3390 92942 3442
rect 97234 3390 97246 3442
rect 97298 3390 97310 3442
rect 100706 3390 100718 3442
rect 100770 3390 100782 3442
rect 101938 3390 101950 3442
rect 102002 3390 102014 3442
rect 104066 3390 104078 3442
rect 104130 3390 104142 3442
rect 106418 3390 106430 3442
rect 106482 3390 106494 3442
rect 108994 3390 109006 3442
rect 109058 3390 109070 3442
rect 111906 3390 111918 3442
rect 111970 3390 111982 3442
rect 116386 3390 116398 3442
rect 116450 3390 116462 3442
rect 120306 3390 120318 3442
rect 120370 3390 120382 3442
rect 5854 3378 5906 3390
rect 121774 3378 121826 3390
rect 130174 3442 130226 3454
rect 130174 3378 130226 3390
rect 133310 3442 133362 3454
rect 133310 3378 133362 3390
rect 135102 3442 135154 3454
rect 135102 3378 135154 3390
rect 136334 3442 136386 3454
rect 136334 3378 136386 3390
rect 142046 3442 142098 3454
rect 142046 3378 142098 3390
rect 145630 3442 145682 3454
rect 145630 3378 145682 3390
rect 145966 3442 146018 3454
rect 145966 3378 146018 3390
rect 148654 3442 148706 3454
rect 148654 3378 148706 3390
rect 152910 3442 152962 3454
rect 152910 3378 152962 3390
rect 155038 3442 155090 3454
rect 155038 3378 155090 3390
rect 157390 3442 157442 3454
rect 157390 3378 157442 3390
rect 159854 3442 159906 3454
rect 159854 3378 159906 3390
rect 162878 3442 162930 3454
rect 162878 3378 162930 3390
rect 164670 3442 164722 3454
rect 164670 3378 164722 3390
rect 166798 3442 166850 3454
rect 166798 3378 166850 3390
rect 168590 3442 168642 3454
rect 168590 3378 168642 3390
rect 171614 3442 171666 3454
rect 171614 3378 171666 3390
rect 14590 3330 14642 3342
rect 14590 3266 14642 3278
rect 25678 3330 25730 3342
rect 25678 3266 25730 3278
rect 28478 3330 28530 3342
rect 28478 3266 28530 3278
rect 29710 3330 29762 3342
rect 29710 3266 29762 3278
rect 65550 3330 65602 3342
rect 65550 3266 65602 3278
rect 98142 3330 98194 3342
rect 98142 3266 98194 3278
rect 122446 3330 122498 3342
rect 122446 3266 122498 3278
rect 123342 3330 123394 3342
rect 123342 3266 123394 3278
rect 124238 3330 124290 3342
rect 124238 3266 124290 3278
rect 125134 3330 125186 3342
rect 125134 3266 125186 3278
rect 126030 3330 126082 3342
rect 126030 3266 126082 3278
rect 127598 3330 127650 3342
rect 127598 3266 127650 3278
rect 128158 3330 128210 3342
rect 128158 3266 128210 3278
rect 129390 3330 129442 3342
rect 129390 3266 129442 3278
rect 130062 3330 130114 3342
rect 130062 3266 130114 3278
rect 131182 3330 131234 3342
rect 131182 3266 131234 3278
rect 132414 3330 132466 3342
rect 132414 3266 132466 3278
rect 132974 3330 133026 3342
rect 132974 3266 133026 3278
rect 133870 3330 133922 3342
rect 133870 3266 133922 3278
rect 135998 3330 136050 3342
rect 135998 3266 136050 3278
rect 136894 3330 136946 3342
rect 136894 3266 136946 3278
rect 137790 3330 137842 3342
rect 137790 3266 137842 3278
rect 139358 3330 139410 3342
rect 139358 3266 139410 3278
rect 139918 3330 139970 3342
rect 139918 3266 139970 3278
rect 140814 3330 140866 3342
rect 140814 3266 140866 3278
rect 141710 3330 141762 3342
rect 141710 3266 141762 3278
rect 142942 3330 142994 3342
rect 142942 3266 142994 3278
rect 143838 3330 143890 3342
rect 143838 3266 143890 3278
rect 144734 3330 144786 3342
rect 144734 3266 144786 3278
rect 146862 3330 146914 3342
rect 146862 3266 146914 3278
rect 147758 3330 147810 3342
rect 147758 3266 147810 3278
rect 149550 3330 149602 3342
rect 149550 3266 149602 3278
rect 150782 3330 150834 3342
rect 150782 3266 150834 3278
rect 151678 3330 151730 3342
rect 151678 3266 151730 3278
rect 152574 3330 152626 3342
rect 152574 3266 152626 3278
rect 153470 3330 153522 3342
rect 153470 3266 153522 3278
rect 154702 3330 154754 3342
rect 154702 3266 154754 3278
rect 155598 3330 155650 3342
rect 155598 3266 155650 3278
rect 156494 3330 156546 3342
rect 156494 3266 156546 3278
rect 158622 3330 158674 3342
rect 158622 3266 158674 3278
rect 159518 3330 159570 3342
rect 159518 3266 159570 3278
rect 160414 3330 160466 3342
rect 160414 3266 160466 3278
rect 161310 3330 161362 3342
rect 161310 3266 161362 3278
rect 162542 3330 162594 3342
rect 162542 3266 162594 3278
rect 163438 3330 163490 3342
rect 163438 3266 163490 3278
rect 164334 3330 164386 3342
rect 164334 3266 164386 3278
rect 165230 3330 165282 3342
rect 165230 3266 165282 3278
rect 166462 3330 166514 3342
rect 166462 3266 166514 3278
rect 167358 3330 167410 3342
rect 167358 3266 167410 3278
rect 168254 3330 168306 3342
rect 168254 3266 168306 3278
rect 169150 3330 169202 3342
rect 169150 3266 169202 3278
rect 170382 3330 170434 3342
rect 170382 3266 170434 3278
rect 171278 3330 171330 3342
rect 171278 3266 171330 3278
rect 172174 3330 172226 3342
rect 172174 3266 172226 3278
rect 173070 3330 173122 3342
rect 173070 3266 173122 3278
rect 174302 3330 174354 3342
rect 174302 3266 174354 3278
rect 174974 3330 175026 3342
rect 174974 3266 175026 3278
rect 1344 3162 178640 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 81278 3162
rect 81330 3110 81382 3162
rect 81434 3110 81486 3162
rect 81538 3110 111998 3162
rect 112050 3110 112102 3162
rect 112154 3110 112206 3162
rect 112258 3110 142718 3162
rect 142770 3110 142822 3162
rect 142874 3110 142926 3162
rect 142978 3110 173438 3162
rect 173490 3110 173542 3162
rect 173594 3110 173646 3162
rect 173698 3110 178640 3162
rect 1344 3076 178640 3110
rect 128706 2942 128718 2994
rect 128770 2991 128782 2994
rect 129378 2991 129390 2994
rect 128770 2945 129390 2991
rect 128770 2942 128782 2945
rect 129378 2942 129390 2945
rect 129442 2942 129454 2994
rect 173394 1710 173406 1762
rect 173458 1759 173470 1762
rect 174290 1759 174302 1762
rect 173458 1713 174302 1759
rect 173458 1710 173470 1713
rect 174290 1710 174302 1713
rect 174354 1710 174366 1762
<< via1 >>
rect 158174 117070 158226 117122
rect 159294 117070 159346 117122
rect 30494 116958 30546 117010
rect 31614 116958 31666 117010
rect 77534 116958 77586 117010
rect 78654 116958 78706 117010
rect 111134 116958 111186 117010
rect 112254 116958 112306 117010
rect 112702 116958 112754 117010
rect 113598 116958 113650 117010
rect 134654 116958 134706 117010
rect 135774 116958 135826 117010
rect 136222 116958 136274 117010
rect 137566 116958 137618 117010
rect 159742 116958 159794 117010
rect 160414 116958 160466 117010
rect 4478 116790 4530 116842
rect 4582 116790 4634 116842
rect 4686 116790 4738 116842
rect 35198 116790 35250 116842
rect 35302 116790 35354 116842
rect 35406 116790 35458 116842
rect 65918 116790 65970 116842
rect 66022 116790 66074 116842
rect 66126 116790 66178 116842
rect 96638 116790 96690 116842
rect 96742 116790 96794 116842
rect 96846 116790 96898 116842
rect 127358 116790 127410 116842
rect 127462 116790 127514 116842
rect 127566 116790 127618 116842
rect 158078 116790 158130 116842
rect 158182 116790 158234 116842
rect 158286 116790 158338 116842
rect 3390 116510 3442 116562
rect 5966 116510 6018 116562
rect 8430 116510 8482 116562
rect 10110 116510 10162 116562
rect 14366 116510 14418 116562
rect 19070 116510 19122 116562
rect 22206 116510 22258 116562
rect 23550 116510 23602 116562
rect 27358 116510 27410 116562
rect 29486 116510 29538 116562
rect 31950 116510 32002 116562
rect 33630 116510 33682 116562
rect 37886 116510 37938 116562
rect 42590 116510 42642 116562
rect 45726 116510 45778 116562
rect 47070 116510 47122 116562
rect 50878 116510 50930 116562
rect 53006 116510 53058 116562
rect 55470 116510 55522 116562
rect 57150 116510 57202 116562
rect 61406 116510 61458 116562
rect 66110 116510 66162 116562
rect 69246 116510 69298 116562
rect 70590 116510 70642 116562
rect 74398 116510 74450 116562
rect 76526 116510 76578 116562
rect 78990 116510 79042 116562
rect 80670 116510 80722 116562
rect 84926 116510 84978 116562
rect 89630 116510 89682 116562
rect 93214 116510 93266 116562
rect 97918 116510 97970 116562
rect 100046 116510 100098 116562
rect 102510 116510 102562 116562
rect 104190 116510 104242 116562
rect 108334 116510 108386 116562
rect 112254 116510 112306 116562
rect 113598 116510 113650 116562
rect 116734 116510 116786 116562
rect 121438 116510 121490 116562
rect 124014 116510 124066 116562
rect 126030 116510 126082 116562
rect 127934 116510 127986 116562
rect 131854 116510 131906 116562
rect 135774 116510 135826 116562
rect 137566 116510 137618 116562
rect 140254 116510 140306 116562
rect 144958 116510 145010 116562
rect 147534 116510 147586 116562
rect 149550 116510 149602 116562
rect 151454 116510 151506 116562
rect 155374 116510 155426 116562
rect 159294 116510 159346 116562
rect 163774 116510 163826 116562
rect 168478 116510 168530 116562
rect 173070 116510 173122 116562
rect 4398 116398 4450 116450
rect 6750 116398 6802 116450
rect 7646 116398 7698 116450
rect 10894 116398 10946 116450
rect 15374 116398 15426 116450
rect 19854 116398 19906 116450
rect 20526 116398 20578 116450
rect 21758 116398 21810 116450
rect 24558 116398 24610 116450
rect 26686 116398 26738 116450
rect 30494 116398 30546 116450
rect 31166 116398 31218 116450
rect 34414 116398 34466 116450
rect 38894 116398 38946 116450
rect 43598 116398 43650 116450
rect 45278 116398 45330 116450
rect 48078 116398 48130 116450
rect 50206 116398 50258 116450
rect 53790 116398 53842 116450
rect 54686 116398 54738 116450
rect 57934 116398 57986 116450
rect 62414 116398 62466 116450
rect 67118 116398 67170 116450
rect 68798 116398 68850 116450
rect 71374 116398 71426 116450
rect 73726 116398 73778 116450
rect 77534 116398 77586 116450
rect 78206 116398 78258 116450
rect 81230 116398 81282 116450
rect 81902 116398 81954 116450
rect 85934 116398 85986 116450
rect 90638 116398 90690 116450
rect 92542 116398 92594 116450
rect 97246 116398 97298 116450
rect 101054 116398 101106 116450
rect 101726 116398 101778 116450
rect 104974 116398 105026 116450
rect 107662 116398 107714 116450
rect 111582 116398 111634 116450
rect 114382 116398 114434 116450
rect 116062 116398 116114 116450
rect 120990 116398 121042 116450
rect 123342 116398 123394 116450
rect 125246 116398 125298 116450
rect 127262 116398 127314 116450
rect 131182 116398 131234 116450
rect 135102 116398 135154 116450
rect 136894 116398 136946 116450
rect 139582 116398 139634 116450
rect 144286 116398 144338 116450
rect 146078 116398 146130 116450
rect 146862 116398 146914 116450
rect 148766 116398 148818 116450
rect 150782 116398 150834 116450
rect 154702 116398 154754 116450
rect 158622 116398 158674 116450
rect 163102 116398 163154 116450
rect 167806 116398 167858 116450
rect 172286 116398 172338 116450
rect 39342 116286 39394 116338
rect 160414 116286 160466 116338
rect 164894 116286 164946 116338
rect 170382 116286 170434 116338
rect 174302 116286 174354 116338
rect 177214 116286 177266 116338
rect 11342 116174 11394 116226
rect 15822 116174 15874 116226
rect 25230 116174 25282 116226
rect 34862 116174 34914 116226
rect 44046 116174 44098 116226
rect 48750 116174 48802 116226
rect 58382 116174 58434 116226
rect 62862 116174 62914 116226
rect 67566 116174 67618 116226
rect 72270 116174 72322 116226
rect 86382 116174 86434 116226
rect 91086 116174 91138 116226
rect 105422 116174 105474 116226
rect 122558 116174 122610 116226
rect 19838 116006 19890 116058
rect 19942 116006 19994 116058
rect 20046 116006 20098 116058
rect 50558 116006 50610 116058
rect 50662 116006 50714 116058
rect 50766 116006 50818 116058
rect 81278 116006 81330 116058
rect 81382 116006 81434 116058
rect 81486 116006 81538 116058
rect 111998 116006 112050 116058
rect 112102 116006 112154 116058
rect 112206 116006 112258 116058
rect 142718 116006 142770 116058
rect 142822 116006 142874 116058
rect 142926 116006 142978 116058
rect 173438 116006 173490 116058
rect 173542 116006 173594 116058
rect 173646 116006 173698 116058
rect 4398 115838 4450 115890
rect 7534 115838 7586 115890
rect 21758 115838 21810 115890
rect 26462 115838 26514 115890
rect 31166 115838 31218 115890
rect 31614 115838 31666 115890
rect 45278 115838 45330 115890
rect 49982 115838 50034 115890
rect 54686 115838 54738 115890
rect 68798 115838 68850 115890
rect 73726 115838 73778 115890
rect 78206 115838 78258 115890
rect 78654 115838 78706 115890
rect 92318 115838 92370 115890
rect 97246 115838 97298 115890
rect 101726 115838 101778 115890
rect 106318 115838 106370 115890
rect 111134 115838 111186 115890
rect 115838 115838 115890 115890
rect 121102 115838 121154 115890
rect 125134 115838 125186 115890
rect 126926 115838 126978 115890
rect 129838 115838 129890 115890
rect 134654 115838 134706 115890
rect 139358 115838 139410 115890
rect 144062 115838 144114 115890
rect 148766 115838 148818 115890
rect 150446 115838 150498 115890
rect 153470 115838 153522 115890
rect 155262 115838 155314 115890
rect 158174 115838 158226 115890
rect 162878 115838 162930 115890
rect 167582 115838 167634 115890
rect 170942 115838 170994 115890
rect 178110 115838 178162 115890
rect 12014 115726 12066 115778
rect 16942 115726 16994 115778
rect 18622 115726 18674 115778
rect 35534 115726 35586 115778
rect 40574 115726 40626 115778
rect 55134 115726 55186 115778
rect 59054 115726 59106 115778
rect 64094 115726 64146 115778
rect 82574 115726 82626 115778
rect 94446 115726 94498 115778
rect 108558 115726 108610 115778
rect 118526 115726 118578 115778
rect 132638 115726 132690 115778
rect 142046 115726 142098 115778
rect 4734 115614 4786 115666
rect 5182 115614 5234 115666
rect 7198 115614 7250 115666
rect 7982 115614 8034 115666
rect 11118 115614 11170 115666
rect 11678 115614 11730 115666
rect 12574 115614 12626 115666
rect 16046 115614 16098 115666
rect 16718 115614 16770 115666
rect 17726 115614 17778 115666
rect 20862 115614 20914 115666
rect 21534 115614 21586 115666
rect 25566 115614 25618 115666
rect 26238 115614 26290 115666
rect 30270 115614 30322 115666
rect 30942 115614 30994 115666
rect 34638 115614 34690 115666
rect 35198 115614 35250 115666
rect 36094 115614 36146 115666
rect 39678 115614 39730 115666
rect 40238 115614 40290 115666
rect 41582 115614 41634 115666
rect 44382 115614 44434 115666
rect 45054 115614 45106 115666
rect 48750 115614 48802 115666
rect 49758 115614 49810 115666
rect 54462 115614 54514 115666
rect 58718 115614 58770 115666
rect 59614 115614 59666 115666
rect 63758 115614 63810 115666
rect 68574 115614 68626 115666
rect 73502 115614 73554 115666
rect 77982 115614 78034 115666
rect 82238 115614 82290 115666
rect 83134 115614 83186 115666
rect 87278 115614 87330 115666
rect 91982 115614 92034 115666
rect 95342 115614 95394 115666
rect 96462 115614 96514 115666
rect 97582 115614 97634 115666
rect 100830 115614 100882 115666
rect 101390 115614 101442 115666
rect 105422 115614 105474 115666
rect 105982 115614 106034 115666
rect 109230 115614 109282 115666
rect 110798 115614 110850 115666
rect 114942 115614 114994 115666
rect 115502 115614 115554 115666
rect 117630 115614 117682 115666
rect 120318 115614 120370 115666
rect 121326 115614 121378 115666
rect 124238 115614 124290 115666
rect 124798 115614 124850 115666
rect 128942 115614 128994 115666
rect 129614 115614 129666 115666
rect 131742 115614 131794 115666
rect 133758 115614 133810 115666
rect 134318 115614 134370 115666
rect 138462 115614 138514 115666
rect 139134 115614 139186 115666
rect 141150 115614 141202 115666
rect 143166 115614 143218 115666
rect 143838 115614 143890 115666
rect 147870 115614 147922 115666
rect 148542 115614 148594 115666
rect 152126 115614 152178 115666
rect 153246 115614 153298 115666
rect 157278 115614 157330 115666
rect 157838 115614 157890 115666
rect 161982 115614 162034 115666
rect 162542 115614 162594 115666
rect 166686 115614 166738 115666
rect 167246 115614 167298 115666
rect 170046 115614 170098 115666
rect 170606 115614 170658 115666
rect 6638 115502 6690 115554
rect 13246 115502 13298 115554
rect 36766 115502 36818 115554
rect 42254 115502 42306 115554
rect 53790 115502 53842 115554
rect 58158 115502 58210 115554
rect 60286 115502 60338 115554
rect 63198 115502 63250 115554
rect 67902 115502 67954 115554
rect 72606 115502 72658 115554
rect 77310 115502 77362 115554
rect 81678 115502 81730 115554
rect 83806 115502 83858 115554
rect 87950 115502 88002 115554
rect 91422 115502 91474 115554
rect 95902 115502 95954 115554
rect 102174 115502 102226 115554
rect 110014 115502 110066 115554
rect 113038 115502 113090 115554
rect 117182 115502 117234 115554
rect 131294 115502 131346 115554
rect 136894 115502 136946 115554
rect 140702 115502 140754 115554
rect 4478 115222 4530 115274
rect 4582 115222 4634 115274
rect 4686 115222 4738 115274
rect 35198 115222 35250 115274
rect 35302 115222 35354 115274
rect 35406 115222 35458 115274
rect 65918 115222 65970 115274
rect 66022 115222 66074 115274
rect 66126 115222 66178 115274
rect 96638 115222 96690 115274
rect 96742 115222 96794 115274
rect 96846 115222 96898 115274
rect 127358 115222 127410 115274
rect 127462 115222 127514 115274
rect 127566 115222 127618 115274
rect 158078 115222 158130 115274
rect 158182 115222 158234 115274
rect 158286 115222 158338 115274
rect 64990 114942 65042 114994
rect 110462 114942 110514 114994
rect 64318 114830 64370 114882
rect 86718 114830 86770 114882
rect 87614 114830 87666 114882
rect 87278 114718 87330 114770
rect 19838 114438 19890 114490
rect 19942 114438 19994 114490
rect 20046 114438 20098 114490
rect 50558 114438 50610 114490
rect 50662 114438 50714 114490
rect 50766 114438 50818 114490
rect 81278 114438 81330 114490
rect 81382 114438 81434 114490
rect 81486 114438 81538 114490
rect 111998 114438 112050 114490
rect 112102 114438 112154 114490
rect 112206 114438 112258 114490
rect 142718 114438 142770 114490
rect 142822 114438 142874 114490
rect 142926 114438 142978 114490
rect 173438 114438 173490 114490
rect 173542 114438 173594 114490
rect 173646 114438 173698 114490
rect 4478 113654 4530 113706
rect 4582 113654 4634 113706
rect 4686 113654 4738 113706
rect 35198 113654 35250 113706
rect 35302 113654 35354 113706
rect 35406 113654 35458 113706
rect 65918 113654 65970 113706
rect 66022 113654 66074 113706
rect 66126 113654 66178 113706
rect 96638 113654 96690 113706
rect 96742 113654 96794 113706
rect 96846 113654 96898 113706
rect 127358 113654 127410 113706
rect 127462 113654 127514 113706
rect 127566 113654 127618 113706
rect 158078 113654 158130 113706
rect 158182 113654 158234 113706
rect 158286 113654 158338 113706
rect 19838 112870 19890 112922
rect 19942 112870 19994 112922
rect 20046 112870 20098 112922
rect 50558 112870 50610 112922
rect 50662 112870 50714 112922
rect 50766 112870 50818 112922
rect 81278 112870 81330 112922
rect 81382 112870 81434 112922
rect 81486 112870 81538 112922
rect 111998 112870 112050 112922
rect 112102 112870 112154 112922
rect 112206 112870 112258 112922
rect 142718 112870 142770 112922
rect 142822 112870 142874 112922
rect 142926 112870 142978 112922
rect 173438 112870 173490 112922
rect 173542 112870 173594 112922
rect 173646 112870 173698 112922
rect 4478 112086 4530 112138
rect 4582 112086 4634 112138
rect 4686 112086 4738 112138
rect 35198 112086 35250 112138
rect 35302 112086 35354 112138
rect 35406 112086 35458 112138
rect 65918 112086 65970 112138
rect 66022 112086 66074 112138
rect 66126 112086 66178 112138
rect 96638 112086 96690 112138
rect 96742 112086 96794 112138
rect 96846 112086 96898 112138
rect 127358 112086 127410 112138
rect 127462 112086 127514 112138
rect 127566 112086 127618 112138
rect 158078 112086 158130 112138
rect 158182 112086 158234 112138
rect 158286 112086 158338 112138
rect 19838 111302 19890 111354
rect 19942 111302 19994 111354
rect 20046 111302 20098 111354
rect 50558 111302 50610 111354
rect 50662 111302 50714 111354
rect 50766 111302 50818 111354
rect 81278 111302 81330 111354
rect 81382 111302 81434 111354
rect 81486 111302 81538 111354
rect 111998 111302 112050 111354
rect 112102 111302 112154 111354
rect 112206 111302 112258 111354
rect 142718 111302 142770 111354
rect 142822 111302 142874 111354
rect 142926 111302 142978 111354
rect 173438 111302 173490 111354
rect 173542 111302 173594 111354
rect 173646 111302 173698 111354
rect 4478 110518 4530 110570
rect 4582 110518 4634 110570
rect 4686 110518 4738 110570
rect 35198 110518 35250 110570
rect 35302 110518 35354 110570
rect 35406 110518 35458 110570
rect 65918 110518 65970 110570
rect 66022 110518 66074 110570
rect 66126 110518 66178 110570
rect 96638 110518 96690 110570
rect 96742 110518 96794 110570
rect 96846 110518 96898 110570
rect 127358 110518 127410 110570
rect 127462 110518 127514 110570
rect 127566 110518 127618 110570
rect 158078 110518 158130 110570
rect 158182 110518 158234 110570
rect 158286 110518 158338 110570
rect 19838 109734 19890 109786
rect 19942 109734 19994 109786
rect 20046 109734 20098 109786
rect 50558 109734 50610 109786
rect 50662 109734 50714 109786
rect 50766 109734 50818 109786
rect 81278 109734 81330 109786
rect 81382 109734 81434 109786
rect 81486 109734 81538 109786
rect 111998 109734 112050 109786
rect 112102 109734 112154 109786
rect 112206 109734 112258 109786
rect 142718 109734 142770 109786
rect 142822 109734 142874 109786
rect 142926 109734 142978 109786
rect 173438 109734 173490 109786
rect 173542 109734 173594 109786
rect 173646 109734 173698 109786
rect 4478 108950 4530 109002
rect 4582 108950 4634 109002
rect 4686 108950 4738 109002
rect 35198 108950 35250 109002
rect 35302 108950 35354 109002
rect 35406 108950 35458 109002
rect 65918 108950 65970 109002
rect 66022 108950 66074 109002
rect 66126 108950 66178 109002
rect 96638 108950 96690 109002
rect 96742 108950 96794 109002
rect 96846 108950 96898 109002
rect 127358 108950 127410 109002
rect 127462 108950 127514 109002
rect 127566 108950 127618 109002
rect 158078 108950 158130 109002
rect 158182 108950 158234 109002
rect 158286 108950 158338 109002
rect 19838 108166 19890 108218
rect 19942 108166 19994 108218
rect 20046 108166 20098 108218
rect 50558 108166 50610 108218
rect 50662 108166 50714 108218
rect 50766 108166 50818 108218
rect 81278 108166 81330 108218
rect 81382 108166 81434 108218
rect 81486 108166 81538 108218
rect 111998 108166 112050 108218
rect 112102 108166 112154 108218
rect 112206 108166 112258 108218
rect 142718 108166 142770 108218
rect 142822 108166 142874 108218
rect 142926 108166 142978 108218
rect 173438 108166 173490 108218
rect 173542 108166 173594 108218
rect 173646 108166 173698 108218
rect 4478 107382 4530 107434
rect 4582 107382 4634 107434
rect 4686 107382 4738 107434
rect 35198 107382 35250 107434
rect 35302 107382 35354 107434
rect 35406 107382 35458 107434
rect 65918 107382 65970 107434
rect 66022 107382 66074 107434
rect 66126 107382 66178 107434
rect 96638 107382 96690 107434
rect 96742 107382 96794 107434
rect 96846 107382 96898 107434
rect 127358 107382 127410 107434
rect 127462 107382 127514 107434
rect 127566 107382 127618 107434
rect 158078 107382 158130 107434
rect 158182 107382 158234 107434
rect 158286 107382 158338 107434
rect 19838 106598 19890 106650
rect 19942 106598 19994 106650
rect 20046 106598 20098 106650
rect 50558 106598 50610 106650
rect 50662 106598 50714 106650
rect 50766 106598 50818 106650
rect 81278 106598 81330 106650
rect 81382 106598 81434 106650
rect 81486 106598 81538 106650
rect 111998 106598 112050 106650
rect 112102 106598 112154 106650
rect 112206 106598 112258 106650
rect 142718 106598 142770 106650
rect 142822 106598 142874 106650
rect 142926 106598 142978 106650
rect 173438 106598 173490 106650
rect 173542 106598 173594 106650
rect 173646 106598 173698 106650
rect 4478 105814 4530 105866
rect 4582 105814 4634 105866
rect 4686 105814 4738 105866
rect 35198 105814 35250 105866
rect 35302 105814 35354 105866
rect 35406 105814 35458 105866
rect 65918 105814 65970 105866
rect 66022 105814 66074 105866
rect 66126 105814 66178 105866
rect 96638 105814 96690 105866
rect 96742 105814 96794 105866
rect 96846 105814 96898 105866
rect 127358 105814 127410 105866
rect 127462 105814 127514 105866
rect 127566 105814 127618 105866
rect 158078 105814 158130 105866
rect 158182 105814 158234 105866
rect 158286 105814 158338 105866
rect 19838 105030 19890 105082
rect 19942 105030 19994 105082
rect 20046 105030 20098 105082
rect 50558 105030 50610 105082
rect 50662 105030 50714 105082
rect 50766 105030 50818 105082
rect 81278 105030 81330 105082
rect 81382 105030 81434 105082
rect 81486 105030 81538 105082
rect 111998 105030 112050 105082
rect 112102 105030 112154 105082
rect 112206 105030 112258 105082
rect 142718 105030 142770 105082
rect 142822 105030 142874 105082
rect 142926 105030 142978 105082
rect 173438 105030 173490 105082
rect 173542 105030 173594 105082
rect 173646 105030 173698 105082
rect 4478 104246 4530 104298
rect 4582 104246 4634 104298
rect 4686 104246 4738 104298
rect 35198 104246 35250 104298
rect 35302 104246 35354 104298
rect 35406 104246 35458 104298
rect 65918 104246 65970 104298
rect 66022 104246 66074 104298
rect 66126 104246 66178 104298
rect 96638 104246 96690 104298
rect 96742 104246 96794 104298
rect 96846 104246 96898 104298
rect 127358 104246 127410 104298
rect 127462 104246 127514 104298
rect 127566 104246 127618 104298
rect 158078 104246 158130 104298
rect 158182 104246 158234 104298
rect 158286 104246 158338 104298
rect 19838 103462 19890 103514
rect 19942 103462 19994 103514
rect 20046 103462 20098 103514
rect 50558 103462 50610 103514
rect 50662 103462 50714 103514
rect 50766 103462 50818 103514
rect 81278 103462 81330 103514
rect 81382 103462 81434 103514
rect 81486 103462 81538 103514
rect 111998 103462 112050 103514
rect 112102 103462 112154 103514
rect 112206 103462 112258 103514
rect 142718 103462 142770 103514
rect 142822 103462 142874 103514
rect 142926 103462 142978 103514
rect 173438 103462 173490 103514
rect 173542 103462 173594 103514
rect 173646 103462 173698 103514
rect 4478 102678 4530 102730
rect 4582 102678 4634 102730
rect 4686 102678 4738 102730
rect 35198 102678 35250 102730
rect 35302 102678 35354 102730
rect 35406 102678 35458 102730
rect 65918 102678 65970 102730
rect 66022 102678 66074 102730
rect 66126 102678 66178 102730
rect 96638 102678 96690 102730
rect 96742 102678 96794 102730
rect 96846 102678 96898 102730
rect 127358 102678 127410 102730
rect 127462 102678 127514 102730
rect 127566 102678 127618 102730
rect 158078 102678 158130 102730
rect 158182 102678 158234 102730
rect 158286 102678 158338 102730
rect 19838 101894 19890 101946
rect 19942 101894 19994 101946
rect 20046 101894 20098 101946
rect 50558 101894 50610 101946
rect 50662 101894 50714 101946
rect 50766 101894 50818 101946
rect 81278 101894 81330 101946
rect 81382 101894 81434 101946
rect 81486 101894 81538 101946
rect 111998 101894 112050 101946
rect 112102 101894 112154 101946
rect 112206 101894 112258 101946
rect 142718 101894 142770 101946
rect 142822 101894 142874 101946
rect 142926 101894 142978 101946
rect 173438 101894 173490 101946
rect 173542 101894 173594 101946
rect 173646 101894 173698 101946
rect 4478 101110 4530 101162
rect 4582 101110 4634 101162
rect 4686 101110 4738 101162
rect 35198 101110 35250 101162
rect 35302 101110 35354 101162
rect 35406 101110 35458 101162
rect 65918 101110 65970 101162
rect 66022 101110 66074 101162
rect 66126 101110 66178 101162
rect 96638 101110 96690 101162
rect 96742 101110 96794 101162
rect 96846 101110 96898 101162
rect 127358 101110 127410 101162
rect 127462 101110 127514 101162
rect 127566 101110 127618 101162
rect 158078 101110 158130 101162
rect 158182 101110 158234 101162
rect 158286 101110 158338 101162
rect 19838 100326 19890 100378
rect 19942 100326 19994 100378
rect 20046 100326 20098 100378
rect 50558 100326 50610 100378
rect 50662 100326 50714 100378
rect 50766 100326 50818 100378
rect 81278 100326 81330 100378
rect 81382 100326 81434 100378
rect 81486 100326 81538 100378
rect 111998 100326 112050 100378
rect 112102 100326 112154 100378
rect 112206 100326 112258 100378
rect 142718 100326 142770 100378
rect 142822 100326 142874 100378
rect 142926 100326 142978 100378
rect 173438 100326 173490 100378
rect 173542 100326 173594 100378
rect 173646 100326 173698 100378
rect 4478 99542 4530 99594
rect 4582 99542 4634 99594
rect 4686 99542 4738 99594
rect 35198 99542 35250 99594
rect 35302 99542 35354 99594
rect 35406 99542 35458 99594
rect 65918 99542 65970 99594
rect 66022 99542 66074 99594
rect 66126 99542 66178 99594
rect 96638 99542 96690 99594
rect 96742 99542 96794 99594
rect 96846 99542 96898 99594
rect 127358 99542 127410 99594
rect 127462 99542 127514 99594
rect 127566 99542 127618 99594
rect 158078 99542 158130 99594
rect 158182 99542 158234 99594
rect 158286 99542 158338 99594
rect 19838 98758 19890 98810
rect 19942 98758 19994 98810
rect 20046 98758 20098 98810
rect 50558 98758 50610 98810
rect 50662 98758 50714 98810
rect 50766 98758 50818 98810
rect 81278 98758 81330 98810
rect 81382 98758 81434 98810
rect 81486 98758 81538 98810
rect 111998 98758 112050 98810
rect 112102 98758 112154 98810
rect 112206 98758 112258 98810
rect 142718 98758 142770 98810
rect 142822 98758 142874 98810
rect 142926 98758 142978 98810
rect 173438 98758 173490 98810
rect 173542 98758 173594 98810
rect 173646 98758 173698 98810
rect 4478 97974 4530 98026
rect 4582 97974 4634 98026
rect 4686 97974 4738 98026
rect 35198 97974 35250 98026
rect 35302 97974 35354 98026
rect 35406 97974 35458 98026
rect 65918 97974 65970 98026
rect 66022 97974 66074 98026
rect 66126 97974 66178 98026
rect 96638 97974 96690 98026
rect 96742 97974 96794 98026
rect 96846 97974 96898 98026
rect 127358 97974 127410 98026
rect 127462 97974 127514 98026
rect 127566 97974 127618 98026
rect 158078 97974 158130 98026
rect 158182 97974 158234 98026
rect 158286 97974 158338 98026
rect 19838 97190 19890 97242
rect 19942 97190 19994 97242
rect 20046 97190 20098 97242
rect 50558 97190 50610 97242
rect 50662 97190 50714 97242
rect 50766 97190 50818 97242
rect 81278 97190 81330 97242
rect 81382 97190 81434 97242
rect 81486 97190 81538 97242
rect 111998 97190 112050 97242
rect 112102 97190 112154 97242
rect 112206 97190 112258 97242
rect 142718 97190 142770 97242
rect 142822 97190 142874 97242
rect 142926 97190 142978 97242
rect 173438 97190 173490 97242
rect 173542 97190 173594 97242
rect 173646 97190 173698 97242
rect 4478 96406 4530 96458
rect 4582 96406 4634 96458
rect 4686 96406 4738 96458
rect 35198 96406 35250 96458
rect 35302 96406 35354 96458
rect 35406 96406 35458 96458
rect 65918 96406 65970 96458
rect 66022 96406 66074 96458
rect 66126 96406 66178 96458
rect 96638 96406 96690 96458
rect 96742 96406 96794 96458
rect 96846 96406 96898 96458
rect 127358 96406 127410 96458
rect 127462 96406 127514 96458
rect 127566 96406 127618 96458
rect 158078 96406 158130 96458
rect 158182 96406 158234 96458
rect 158286 96406 158338 96458
rect 19838 95622 19890 95674
rect 19942 95622 19994 95674
rect 20046 95622 20098 95674
rect 50558 95622 50610 95674
rect 50662 95622 50714 95674
rect 50766 95622 50818 95674
rect 81278 95622 81330 95674
rect 81382 95622 81434 95674
rect 81486 95622 81538 95674
rect 111998 95622 112050 95674
rect 112102 95622 112154 95674
rect 112206 95622 112258 95674
rect 142718 95622 142770 95674
rect 142822 95622 142874 95674
rect 142926 95622 142978 95674
rect 173438 95622 173490 95674
rect 173542 95622 173594 95674
rect 173646 95622 173698 95674
rect 4478 94838 4530 94890
rect 4582 94838 4634 94890
rect 4686 94838 4738 94890
rect 35198 94838 35250 94890
rect 35302 94838 35354 94890
rect 35406 94838 35458 94890
rect 65918 94838 65970 94890
rect 66022 94838 66074 94890
rect 66126 94838 66178 94890
rect 96638 94838 96690 94890
rect 96742 94838 96794 94890
rect 96846 94838 96898 94890
rect 127358 94838 127410 94890
rect 127462 94838 127514 94890
rect 127566 94838 127618 94890
rect 158078 94838 158130 94890
rect 158182 94838 158234 94890
rect 158286 94838 158338 94890
rect 19838 94054 19890 94106
rect 19942 94054 19994 94106
rect 20046 94054 20098 94106
rect 50558 94054 50610 94106
rect 50662 94054 50714 94106
rect 50766 94054 50818 94106
rect 81278 94054 81330 94106
rect 81382 94054 81434 94106
rect 81486 94054 81538 94106
rect 111998 94054 112050 94106
rect 112102 94054 112154 94106
rect 112206 94054 112258 94106
rect 142718 94054 142770 94106
rect 142822 94054 142874 94106
rect 142926 94054 142978 94106
rect 173438 94054 173490 94106
rect 173542 94054 173594 94106
rect 173646 94054 173698 94106
rect 4478 93270 4530 93322
rect 4582 93270 4634 93322
rect 4686 93270 4738 93322
rect 35198 93270 35250 93322
rect 35302 93270 35354 93322
rect 35406 93270 35458 93322
rect 65918 93270 65970 93322
rect 66022 93270 66074 93322
rect 66126 93270 66178 93322
rect 96638 93270 96690 93322
rect 96742 93270 96794 93322
rect 96846 93270 96898 93322
rect 127358 93270 127410 93322
rect 127462 93270 127514 93322
rect 127566 93270 127618 93322
rect 158078 93270 158130 93322
rect 158182 93270 158234 93322
rect 158286 93270 158338 93322
rect 19838 92486 19890 92538
rect 19942 92486 19994 92538
rect 20046 92486 20098 92538
rect 50558 92486 50610 92538
rect 50662 92486 50714 92538
rect 50766 92486 50818 92538
rect 81278 92486 81330 92538
rect 81382 92486 81434 92538
rect 81486 92486 81538 92538
rect 111998 92486 112050 92538
rect 112102 92486 112154 92538
rect 112206 92486 112258 92538
rect 142718 92486 142770 92538
rect 142822 92486 142874 92538
rect 142926 92486 142978 92538
rect 173438 92486 173490 92538
rect 173542 92486 173594 92538
rect 173646 92486 173698 92538
rect 4478 91702 4530 91754
rect 4582 91702 4634 91754
rect 4686 91702 4738 91754
rect 35198 91702 35250 91754
rect 35302 91702 35354 91754
rect 35406 91702 35458 91754
rect 65918 91702 65970 91754
rect 66022 91702 66074 91754
rect 66126 91702 66178 91754
rect 96638 91702 96690 91754
rect 96742 91702 96794 91754
rect 96846 91702 96898 91754
rect 127358 91702 127410 91754
rect 127462 91702 127514 91754
rect 127566 91702 127618 91754
rect 158078 91702 158130 91754
rect 158182 91702 158234 91754
rect 158286 91702 158338 91754
rect 19838 90918 19890 90970
rect 19942 90918 19994 90970
rect 20046 90918 20098 90970
rect 50558 90918 50610 90970
rect 50662 90918 50714 90970
rect 50766 90918 50818 90970
rect 81278 90918 81330 90970
rect 81382 90918 81434 90970
rect 81486 90918 81538 90970
rect 111998 90918 112050 90970
rect 112102 90918 112154 90970
rect 112206 90918 112258 90970
rect 142718 90918 142770 90970
rect 142822 90918 142874 90970
rect 142926 90918 142978 90970
rect 173438 90918 173490 90970
rect 173542 90918 173594 90970
rect 173646 90918 173698 90970
rect 4478 90134 4530 90186
rect 4582 90134 4634 90186
rect 4686 90134 4738 90186
rect 35198 90134 35250 90186
rect 35302 90134 35354 90186
rect 35406 90134 35458 90186
rect 65918 90134 65970 90186
rect 66022 90134 66074 90186
rect 66126 90134 66178 90186
rect 96638 90134 96690 90186
rect 96742 90134 96794 90186
rect 96846 90134 96898 90186
rect 127358 90134 127410 90186
rect 127462 90134 127514 90186
rect 127566 90134 127618 90186
rect 158078 90134 158130 90186
rect 158182 90134 158234 90186
rect 158286 90134 158338 90186
rect 19838 89350 19890 89402
rect 19942 89350 19994 89402
rect 20046 89350 20098 89402
rect 50558 89350 50610 89402
rect 50662 89350 50714 89402
rect 50766 89350 50818 89402
rect 81278 89350 81330 89402
rect 81382 89350 81434 89402
rect 81486 89350 81538 89402
rect 111998 89350 112050 89402
rect 112102 89350 112154 89402
rect 112206 89350 112258 89402
rect 142718 89350 142770 89402
rect 142822 89350 142874 89402
rect 142926 89350 142978 89402
rect 173438 89350 173490 89402
rect 173542 89350 173594 89402
rect 173646 89350 173698 89402
rect 4478 88566 4530 88618
rect 4582 88566 4634 88618
rect 4686 88566 4738 88618
rect 35198 88566 35250 88618
rect 35302 88566 35354 88618
rect 35406 88566 35458 88618
rect 65918 88566 65970 88618
rect 66022 88566 66074 88618
rect 66126 88566 66178 88618
rect 96638 88566 96690 88618
rect 96742 88566 96794 88618
rect 96846 88566 96898 88618
rect 127358 88566 127410 88618
rect 127462 88566 127514 88618
rect 127566 88566 127618 88618
rect 158078 88566 158130 88618
rect 158182 88566 158234 88618
rect 158286 88566 158338 88618
rect 19838 87782 19890 87834
rect 19942 87782 19994 87834
rect 20046 87782 20098 87834
rect 50558 87782 50610 87834
rect 50662 87782 50714 87834
rect 50766 87782 50818 87834
rect 81278 87782 81330 87834
rect 81382 87782 81434 87834
rect 81486 87782 81538 87834
rect 111998 87782 112050 87834
rect 112102 87782 112154 87834
rect 112206 87782 112258 87834
rect 142718 87782 142770 87834
rect 142822 87782 142874 87834
rect 142926 87782 142978 87834
rect 173438 87782 173490 87834
rect 173542 87782 173594 87834
rect 173646 87782 173698 87834
rect 4478 86998 4530 87050
rect 4582 86998 4634 87050
rect 4686 86998 4738 87050
rect 35198 86998 35250 87050
rect 35302 86998 35354 87050
rect 35406 86998 35458 87050
rect 65918 86998 65970 87050
rect 66022 86998 66074 87050
rect 66126 86998 66178 87050
rect 96638 86998 96690 87050
rect 96742 86998 96794 87050
rect 96846 86998 96898 87050
rect 127358 86998 127410 87050
rect 127462 86998 127514 87050
rect 127566 86998 127618 87050
rect 158078 86998 158130 87050
rect 158182 86998 158234 87050
rect 158286 86998 158338 87050
rect 19838 86214 19890 86266
rect 19942 86214 19994 86266
rect 20046 86214 20098 86266
rect 50558 86214 50610 86266
rect 50662 86214 50714 86266
rect 50766 86214 50818 86266
rect 81278 86214 81330 86266
rect 81382 86214 81434 86266
rect 81486 86214 81538 86266
rect 111998 86214 112050 86266
rect 112102 86214 112154 86266
rect 112206 86214 112258 86266
rect 142718 86214 142770 86266
rect 142822 86214 142874 86266
rect 142926 86214 142978 86266
rect 173438 86214 173490 86266
rect 173542 86214 173594 86266
rect 173646 86214 173698 86266
rect 4478 85430 4530 85482
rect 4582 85430 4634 85482
rect 4686 85430 4738 85482
rect 35198 85430 35250 85482
rect 35302 85430 35354 85482
rect 35406 85430 35458 85482
rect 65918 85430 65970 85482
rect 66022 85430 66074 85482
rect 66126 85430 66178 85482
rect 96638 85430 96690 85482
rect 96742 85430 96794 85482
rect 96846 85430 96898 85482
rect 127358 85430 127410 85482
rect 127462 85430 127514 85482
rect 127566 85430 127618 85482
rect 158078 85430 158130 85482
rect 158182 85430 158234 85482
rect 158286 85430 158338 85482
rect 19838 84646 19890 84698
rect 19942 84646 19994 84698
rect 20046 84646 20098 84698
rect 50558 84646 50610 84698
rect 50662 84646 50714 84698
rect 50766 84646 50818 84698
rect 81278 84646 81330 84698
rect 81382 84646 81434 84698
rect 81486 84646 81538 84698
rect 111998 84646 112050 84698
rect 112102 84646 112154 84698
rect 112206 84646 112258 84698
rect 142718 84646 142770 84698
rect 142822 84646 142874 84698
rect 142926 84646 142978 84698
rect 173438 84646 173490 84698
rect 173542 84646 173594 84698
rect 173646 84646 173698 84698
rect 4478 83862 4530 83914
rect 4582 83862 4634 83914
rect 4686 83862 4738 83914
rect 35198 83862 35250 83914
rect 35302 83862 35354 83914
rect 35406 83862 35458 83914
rect 65918 83862 65970 83914
rect 66022 83862 66074 83914
rect 66126 83862 66178 83914
rect 96638 83862 96690 83914
rect 96742 83862 96794 83914
rect 96846 83862 96898 83914
rect 127358 83862 127410 83914
rect 127462 83862 127514 83914
rect 127566 83862 127618 83914
rect 158078 83862 158130 83914
rect 158182 83862 158234 83914
rect 158286 83862 158338 83914
rect 19838 83078 19890 83130
rect 19942 83078 19994 83130
rect 20046 83078 20098 83130
rect 50558 83078 50610 83130
rect 50662 83078 50714 83130
rect 50766 83078 50818 83130
rect 81278 83078 81330 83130
rect 81382 83078 81434 83130
rect 81486 83078 81538 83130
rect 111998 83078 112050 83130
rect 112102 83078 112154 83130
rect 112206 83078 112258 83130
rect 142718 83078 142770 83130
rect 142822 83078 142874 83130
rect 142926 83078 142978 83130
rect 173438 83078 173490 83130
rect 173542 83078 173594 83130
rect 173646 83078 173698 83130
rect 4478 82294 4530 82346
rect 4582 82294 4634 82346
rect 4686 82294 4738 82346
rect 35198 82294 35250 82346
rect 35302 82294 35354 82346
rect 35406 82294 35458 82346
rect 65918 82294 65970 82346
rect 66022 82294 66074 82346
rect 66126 82294 66178 82346
rect 96638 82294 96690 82346
rect 96742 82294 96794 82346
rect 96846 82294 96898 82346
rect 127358 82294 127410 82346
rect 127462 82294 127514 82346
rect 127566 82294 127618 82346
rect 158078 82294 158130 82346
rect 158182 82294 158234 82346
rect 158286 82294 158338 82346
rect 19838 81510 19890 81562
rect 19942 81510 19994 81562
rect 20046 81510 20098 81562
rect 50558 81510 50610 81562
rect 50662 81510 50714 81562
rect 50766 81510 50818 81562
rect 81278 81510 81330 81562
rect 81382 81510 81434 81562
rect 81486 81510 81538 81562
rect 111998 81510 112050 81562
rect 112102 81510 112154 81562
rect 112206 81510 112258 81562
rect 142718 81510 142770 81562
rect 142822 81510 142874 81562
rect 142926 81510 142978 81562
rect 173438 81510 173490 81562
rect 173542 81510 173594 81562
rect 173646 81510 173698 81562
rect 4478 80726 4530 80778
rect 4582 80726 4634 80778
rect 4686 80726 4738 80778
rect 35198 80726 35250 80778
rect 35302 80726 35354 80778
rect 35406 80726 35458 80778
rect 65918 80726 65970 80778
rect 66022 80726 66074 80778
rect 66126 80726 66178 80778
rect 96638 80726 96690 80778
rect 96742 80726 96794 80778
rect 96846 80726 96898 80778
rect 127358 80726 127410 80778
rect 127462 80726 127514 80778
rect 127566 80726 127618 80778
rect 158078 80726 158130 80778
rect 158182 80726 158234 80778
rect 158286 80726 158338 80778
rect 19838 79942 19890 79994
rect 19942 79942 19994 79994
rect 20046 79942 20098 79994
rect 50558 79942 50610 79994
rect 50662 79942 50714 79994
rect 50766 79942 50818 79994
rect 81278 79942 81330 79994
rect 81382 79942 81434 79994
rect 81486 79942 81538 79994
rect 111998 79942 112050 79994
rect 112102 79942 112154 79994
rect 112206 79942 112258 79994
rect 142718 79942 142770 79994
rect 142822 79942 142874 79994
rect 142926 79942 142978 79994
rect 173438 79942 173490 79994
rect 173542 79942 173594 79994
rect 173646 79942 173698 79994
rect 4478 79158 4530 79210
rect 4582 79158 4634 79210
rect 4686 79158 4738 79210
rect 35198 79158 35250 79210
rect 35302 79158 35354 79210
rect 35406 79158 35458 79210
rect 65918 79158 65970 79210
rect 66022 79158 66074 79210
rect 66126 79158 66178 79210
rect 96638 79158 96690 79210
rect 96742 79158 96794 79210
rect 96846 79158 96898 79210
rect 127358 79158 127410 79210
rect 127462 79158 127514 79210
rect 127566 79158 127618 79210
rect 158078 79158 158130 79210
rect 158182 79158 158234 79210
rect 158286 79158 158338 79210
rect 19838 78374 19890 78426
rect 19942 78374 19994 78426
rect 20046 78374 20098 78426
rect 50558 78374 50610 78426
rect 50662 78374 50714 78426
rect 50766 78374 50818 78426
rect 81278 78374 81330 78426
rect 81382 78374 81434 78426
rect 81486 78374 81538 78426
rect 111998 78374 112050 78426
rect 112102 78374 112154 78426
rect 112206 78374 112258 78426
rect 142718 78374 142770 78426
rect 142822 78374 142874 78426
rect 142926 78374 142978 78426
rect 173438 78374 173490 78426
rect 173542 78374 173594 78426
rect 173646 78374 173698 78426
rect 4478 77590 4530 77642
rect 4582 77590 4634 77642
rect 4686 77590 4738 77642
rect 35198 77590 35250 77642
rect 35302 77590 35354 77642
rect 35406 77590 35458 77642
rect 65918 77590 65970 77642
rect 66022 77590 66074 77642
rect 66126 77590 66178 77642
rect 96638 77590 96690 77642
rect 96742 77590 96794 77642
rect 96846 77590 96898 77642
rect 127358 77590 127410 77642
rect 127462 77590 127514 77642
rect 127566 77590 127618 77642
rect 158078 77590 158130 77642
rect 158182 77590 158234 77642
rect 158286 77590 158338 77642
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 81278 76806 81330 76858
rect 81382 76806 81434 76858
rect 81486 76806 81538 76858
rect 111998 76806 112050 76858
rect 112102 76806 112154 76858
rect 112206 76806 112258 76858
rect 142718 76806 142770 76858
rect 142822 76806 142874 76858
rect 142926 76806 142978 76858
rect 173438 76806 173490 76858
rect 173542 76806 173594 76858
rect 173646 76806 173698 76858
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 96638 76022 96690 76074
rect 96742 76022 96794 76074
rect 96846 76022 96898 76074
rect 127358 76022 127410 76074
rect 127462 76022 127514 76074
rect 127566 76022 127618 76074
rect 158078 76022 158130 76074
rect 158182 76022 158234 76074
rect 158286 76022 158338 76074
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 81278 75238 81330 75290
rect 81382 75238 81434 75290
rect 81486 75238 81538 75290
rect 111998 75238 112050 75290
rect 112102 75238 112154 75290
rect 112206 75238 112258 75290
rect 142718 75238 142770 75290
rect 142822 75238 142874 75290
rect 142926 75238 142978 75290
rect 173438 75238 173490 75290
rect 173542 75238 173594 75290
rect 173646 75238 173698 75290
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 96638 74454 96690 74506
rect 96742 74454 96794 74506
rect 96846 74454 96898 74506
rect 127358 74454 127410 74506
rect 127462 74454 127514 74506
rect 127566 74454 127618 74506
rect 158078 74454 158130 74506
rect 158182 74454 158234 74506
rect 158286 74454 158338 74506
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 81278 73670 81330 73722
rect 81382 73670 81434 73722
rect 81486 73670 81538 73722
rect 111998 73670 112050 73722
rect 112102 73670 112154 73722
rect 112206 73670 112258 73722
rect 142718 73670 142770 73722
rect 142822 73670 142874 73722
rect 142926 73670 142978 73722
rect 173438 73670 173490 73722
rect 173542 73670 173594 73722
rect 173646 73670 173698 73722
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 96638 72886 96690 72938
rect 96742 72886 96794 72938
rect 96846 72886 96898 72938
rect 127358 72886 127410 72938
rect 127462 72886 127514 72938
rect 127566 72886 127618 72938
rect 158078 72886 158130 72938
rect 158182 72886 158234 72938
rect 158286 72886 158338 72938
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 81278 72102 81330 72154
rect 81382 72102 81434 72154
rect 81486 72102 81538 72154
rect 111998 72102 112050 72154
rect 112102 72102 112154 72154
rect 112206 72102 112258 72154
rect 142718 72102 142770 72154
rect 142822 72102 142874 72154
rect 142926 72102 142978 72154
rect 173438 72102 173490 72154
rect 173542 72102 173594 72154
rect 173646 72102 173698 72154
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 96638 71318 96690 71370
rect 96742 71318 96794 71370
rect 96846 71318 96898 71370
rect 127358 71318 127410 71370
rect 127462 71318 127514 71370
rect 127566 71318 127618 71370
rect 158078 71318 158130 71370
rect 158182 71318 158234 71370
rect 158286 71318 158338 71370
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 81278 70534 81330 70586
rect 81382 70534 81434 70586
rect 81486 70534 81538 70586
rect 111998 70534 112050 70586
rect 112102 70534 112154 70586
rect 112206 70534 112258 70586
rect 142718 70534 142770 70586
rect 142822 70534 142874 70586
rect 142926 70534 142978 70586
rect 173438 70534 173490 70586
rect 173542 70534 173594 70586
rect 173646 70534 173698 70586
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 96638 69750 96690 69802
rect 96742 69750 96794 69802
rect 96846 69750 96898 69802
rect 127358 69750 127410 69802
rect 127462 69750 127514 69802
rect 127566 69750 127618 69802
rect 158078 69750 158130 69802
rect 158182 69750 158234 69802
rect 158286 69750 158338 69802
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 81278 68966 81330 69018
rect 81382 68966 81434 69018
rect 81486 68966 81538 69018
rect 111998 68966 112050 69018
rect 112102 68966 112154 69018
rect 112206 68966 112258 69018
rect 142718 68966 142770 69018
rect 142822 68966 142874 69018
rect 142926 68966 142978 69018
rect 173438 68966 173490 69018
rect 173542 68966 173594 69018
rect 173646 68966 173698 69018
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 96638 68182 96690 68234
rect 96742 68182 96794 68234
rect 96846 68182 96898 68234
rect 127358 68182 127410 68234
rect 127462 68182 127514 68234
rect 127566 68182 127618 68234
rect 158078 68182 158130 68234
rect 158182 68182 158234 68234
rect 158286 68182 158338 68234
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 81278 67398 81330 67450
rect 81382 67398 81434 67450
rect 81486 67398 81538 67450
rect 111998 67398 112050 67450
rect 112102 67398 112154 67450
rect 112206 67398 112258 67450
rect 142718 67398 142770 67450
rect 142822 67398 142874 67450
rect 142926 67398 142978 67450
rect 173438 67398 173490 67450
rect 173542 67398 173594 67450
rect 173646 67398 173698 67450
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 96638 66614 96690 66666
rect 96742 66614 96794 66666
rect 96846 66614 96898 66666
rect 127358 66614 127410 66666
rect 127462 66614 127514 66666
rect 127566 66614 127618 66666
rect 158078 66614 158130 66666
rect 158182 66614 158234 66666
rect 158286 66614 158338 66666
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 81278 65830 81330 65882
rect 81382 65830 81434 65882
rect 81486 65830 81538 65882
rect 111998 65830 112050 65882
rect 112102 65830 112154 65882
rect 112206 65830 112258 65882
rect 142718 65830 142770 65882
rect 142822 65830 142874 65882
rect 142926 65830 142978 65882
rect 173438 65830 173490 65882
rect 173542 65830 173594 65882
rect 173646 65830 173698 65882
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 96638 65046 96690 65098
rect 96742 65046 96794 65098
rect 96846 65046 96898 65098
rect 127358 65046 127410 65098
rect 127462 65046 127514 65098
rect 127566 65046 127618 65098
rect 158078 65046 158130 65098
rect 158182 65046 158234 65098
rect 158286 65046 158338 65098
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 81278 64262 81330 64314
rect 81382 64262 81434 64314
rect 81486 64262 81538 64314
rect 111998 64262 112050 64314
rect 112102 64262 112154 64314
rect 112206 64262 112258 64314
rect 142718 64262 142770 64314
rect 142822 64262 142874 64314
rect 142926 64262 142978 64314
rect 173438 64262 173490 64314
rect 173542 64262 173594 64314
rect 173646 64262 173698 64314
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 96638 63478 96690 63530
rect 96742 63478 96794 63530
rect 96846 63478 96898 63530
rect 127358 63478 127410 63530
rect 127462 63478 127514 63530
rect 127566 63478 127618 63530
rect 158078 63478 158130 63530
rect 158182 63478 158234 63530
rect 158286 63478 158338 63530
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 81278 62694 81330 62746
rect 81382 62694 81434 62746
rect 81486 62694 81538 62746
rect 111998 62694 112050 62746
rect 112102 62694 112154 62746
rect 112206 62694 112258 62746
rect 142718 62694 142770 62746
rect 142822 62694 142874 62746
rect 142926 62694 142978 62746
rect 173438 62694 173490 62746
rect 173542 62694 173594 62746
rect 173646 62694 173698 62746
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 96638 61910 96690 61962
rect 96742 61910 96794 61962
rect 96846 61910 96898 61962
rect 127358 61910 127410 61962
rect 127462 61910 127514 61962
rect 127566 61910 127618 61962
rect 158078 61910 158130 61962
rect 158182 61910 158234 61962
rect 158286 61910 158338 61962
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 81278 61126 81330 61178
rect 81382 61126 81434 61178
rect 81486 61126 81538 61178
rect 111998 61126 112050 61178
rect 112102 61126 112154 61178
rect 112206 61126 112258 61178
rect 142718 61126 142770 61178
rect 142822 61126 142874 61178
rect 142926 61126 142978 61178
rect 173438 61126 173490 61178
rect 173542 61126 173594 61178
rect 173646 61126 173698 61178
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 96638 60342 96690 60394
rect 96742 60342 96794 60394
rect 96846 60342 96898 60394
rect 127358 60342 127410 60394
rect 127462 60342 127514 60394
rect 127566 60342 127618 60394
rect 158078 60342 158130 60394
rect 158182 60342 158234 60394
rect 158286 60342 158338 60394
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 81278 59558 81330 59610
rect 81382 59558 81434 59610
rect 81486 59558 81538 59610
rect 111998 59558 112050 59610
rect 112102 59558 112154 59610
rect 112206 59558 112258 59610
rect 142718 59558 142770 59610
rect 142822 59558 142874 59610
rect 142926 59558 142978 59610
rect 173438 59558 173490 59610
rect 173542 59558 173594 59610
rect 173646 59558 173698 59610
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 96638 58774 96690 58826
rect 96742 58774 96794 58826
rect 96846 58774 96898 58826
rect 127358 58774 127410 58826
rect 127462 58774 127514 58826
rect 127566 58774 127618 58826
rect 158078 58774 158130 58826
rect 158182 58774 158234 58826
rect 158286 58774 158338 58826
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 81278 57990 81330 58042
rect 81382 57990 81434 58042
rect 81486 57990 81538 58042
rect 111998 57990 112050 58042
rect 112102 57990 112154 58042
rect 112206 57990 112258 58042
rect 142718 57990 142770 58042
rect 142822 57990 142874 58042
rect 142926 57990 142978 58042
rect 173438 57990 173490 58042
rect 173542 57990 173594 58042
rect 173646 57990 173698 58042
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 96638 57206 96690 57258
rect 96742 57206 96794 57258
rect 96846 57206 96898 57258
rect 127358 57206 127410 57258
rect 127462 57206 127514 57258
rect 127566 57206 127618 57258
rect 158078 57206 158130 57258
rect 158182 57206 158234 57258
rect 158286 57206 158338 57258
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 81278 56422 81330 56474
rect 81382 56422 81434 56474
rect 81486 56422 81538 56474
rect 111998 56422 112050 56474
rect 112102 56422 112154 56474
rect 112206 56422 112258 56474
rect 142718 56422 142770 56474
rect 142822 56422 142874 56474
rect 142926 56422 142978 56474
rect 173438 56422 173490 56474
rect 173542 56422 173594 56474
rect 173646 56422 173698 56474
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 96638 55638 96690 55690
rect 96742 55638 96794 55690
rect 96846 55638 96898 55690
rect 127358 55638 127410 55690
rect 127462 55638 127514 55690
rect 127566 55638 127618 55690
rect 158078 55638 158130 55690
rect 158182 55638 158234 55690
rect 158286 55638 158338 55690
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 81278 54854 81330 54906
rect 81382 54854 81434 54906
rect 81486 54854 81538 54906
rect 111998 54854 112050 54906
rect 112102 54854 112154 54906
rect 112206 54854 112258 54906
rect 142718 54854 142770 54906
rect 142822 54854 142874 54906
rect 142926 54854 142978 54906
rect 173438 54854 173490 54906
rect 173542 54854 173594 54906
rect 173646 54854 173698 54906
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 96638 54070 96690 54122
rect 96742 54070 96794 54122
rect 96846 54070 96898 54122
rect 127358 54070 127410 54122
rect 127462 54070 127514 54122
rect 127566 54070 127618 54122
rect 158078 54070 158130 54122
rect 158182 54070 158234 54122
rect 158286 54070 158338 54122
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 81278 53286 81330 53338
rect 81382 53286 81434 53338
rect 81486 53286 81538 53338
rect 111998 53286 112050 53338
rect 112102 53286 112154 53338
rect 112206 53286 112258 53338
rect 142718 53286 142770 53338
rect 142822 53286 142874 53338
rect 142926 53286 142978 53338
rect 173438 53286 173490 53338
rect 173542 53286 173594 53338
rect 173646 53286 173698 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 96638 52502 96690 52554
rect 96742 52502 96794 52554
rect 96846 52502 96898 52554
rect 127358 52502 127410 52554
rect 127462 52502 127514 52554
rect 127566 52502 127618 52554
rect 158078 52502 158130 52554
rect 158182 52502 158234 52554
rect 158286 52502 158338 52554
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 81278 51718 81330 51770
rect 81382 51718 81434 51770
rect 81486 51718 81538 51770
rect 111998 51718 112050 51770
rect 112102 51718 112154 51770
rect 112206 51718 112258 51770
rect 142718 51718 142770 51770
rect 142822 51718 142874 51770
rect 142926 51718 142978 51770
rect 173438 51718 173490 51770
rect 173542 51718 173594 51770
rect 173646 51718 173698 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 96638 50934 96690 50986
rect 96742 50934 96794 50986
rect 96846 50934 96898 50986
rect 127358 50934 127410 50986
rect 127462 50934 127514 50986
rect 127566 50934 127618 50986
rect 158078 50934 158130 50986
rect 158182 50934 158234 50986
rect 158286 50934 158338 50986
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 81278 50150 81330 50202
rect 81382 50150 81434 50202
rect 81486 50150 81538 50202
rect 111998 50150 112050 50202
rect 112102 50150 112154 50202
rect 112206 50150 112258 50202
rect 142718 50150 142770 50202
rect 142822 50150 142874 50202
rect 142926 50150 142978 50202
rect 173438 50150 173490 50202
rect 173542 50150 173594 50202
rect 173646 50150 173698 50202
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 96638 49366 96690 49418
rect 96742 49366 96794 49418
rect 96846 49366 96898 49418
rect 127358 49366 127410 49418
rect 127462 49366 127514 49418
rect 127566 49366 127618 49418
rect 158078 49366 158130 49418
rect 158182 49366 158234 49418
rect 158286 49366 158338 49418
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 81278 48582 81330 48634
rect 81382 48582 81434 48634
rect 81486 48582 81538 48634
rect 111998 48582 112050 48634
rect 112102 48582 112154 48634
rect 112206 48582 112258 48634
rect 142718 48582 142770 48634
rect 142822 48582 142874 48634
rect 142926 48582 142978 48634
rect 173438 48582 173490 48634
rect 173542 48582 173594 48634
rect 173646 48582 173698 48634
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 96638 47798 96690 47850
rect 96742 47798 96794 47850
rect 96846 47798 96898 47850
rect 127358 47798 127410 47850
rect 127462 47798 127514 47850
rect 127566 47798 127618 47850
rect 158078 47798 158130 47850
rect 158182 47798 158234 47850
rect 158286 47798 158338 47850
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 81278 47014 81330 47066
rect 81382 47014 81434 47066
rect 81486 47014 81538 47066
rect 111998 47014 112050 47066
rect 112102 47014 112154 47066
rect 112206 47014 112258 47066
rect 142718 47014 142770 47066
rect 142822 47014 142874 47066
rect 142926 47014 142978 47066
rect 173438 47014 173490 47066
rect 173542 47014 173594 47066
rect 173646 47014 173698 47066
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 96638 46230 96690 46282
rect 96742 46230 96794 46282
rect 96846 46230 96898 46282
rect 127358 46230 127410 46282
rect 127462 46230 127514 46282
rect 127566 46230 127618 46282
rect 158078 46230 158130 46282
rect 158182 46230 158234 46282
rect 158286 46230 158338 46282
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 81278 45446 81330 45498
rect 81382 45446 81434 45498
rect 81486 45446 81538 45498
rect 111998 45446 112050 45498
rect 112102 45446 112154 45498
rect 112206 45446 112258 45498
rect 142718 45446 142770 45498
rect 142822 45446 142874 45498
rect 142926 45446 142978 45498
rect 173438 45446 173490 45498
rect 173542 45446 173594 45498
rect 173646 45446 173698 45498
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 96638 44662 96690 44714
rect 96742 44662 96794 44714
rect 96846 44662 96898 44714
rect 127358 44662 127410 44714
rect 127462 44662 127514 44714
rect 127566 44662 127618 44714
rect 158078 44662 158130 44714
rect 158182 44662 158234 44714
rect 158286 44662 158338 44714
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 81278 43878 81330 43930
rect 81382 43878 81434 43930
rect 81486 43878 81538 43930
rect 111998 43878 112050 43930
rect 112102 43878 112154 43930
rect 112206 43878 112258 43930
rect 142718 43878 142770 43930
rect 142822 43878 142874 43930
rect 142926 43878 142978 43930
rect 173438 43878 173490 43930
rect 173542 43878 173594 43930
rect 173646 43878 173698 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 96638 43094 96690 43146
rect 96742 43094 96794 43146
rect 96846 43094 96898 43146
rect 127358 43094 127410 43146
rect 127462 43094 127514 43146
rect 127566 43094 127618 43146
rect 158078 43094 158130 43146
rect 158182 43094 158234 43146
rect 158286 43094 158338 43146
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 81278 42310 81330 42362
rect 81382 42310 81434 42362
rect 81486 42310 81538 42362
rect 111998 42310 112050 42362
rect 112102 42310 112154 42362
rect 112206 42310 112258 42362
rect 142718 42310 142770 42362
rect 142822 42310 142874 42362
rect 142926 42310 142978 42362
rect 173438 42310 173490 42362
rect 173542 42310 173594 42362
rect 173646 42310 173698 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 96638 41526 96690 41578
rect 96742 41526 96794 41578
rect 96846 41526 96898 41578
rect 127358 41526 127410 41578
rect 127462 41526 127514 41578
rect 127566 41526 127618 41578
rect 158078 41526 158130 41578
rect 158182 41526 158234 41578
rect 158286 41526 158338 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 81278 40742 81330 40794
rect 81382 40742 81434 40794
rect 81486 40742 81538 40794
rect 111998 40742 112050 40794
rect 112102 40742 112154 40794
rect 112206 40742 112258 40794
rect 142718 40742 142770 40794
rect 142822 40742 142874 40794
rect 142926 40742 142978 40794
rect 173438 40742 173490 40794
rect 173542 40742 173594 40794
rect 173646 40742 173698 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 96638 39958 96690 40010
rect 96742 39958 96794 40010
rect 96846 39958 96898 40010
rect 127358 39958 127410 40010
rect 127462 39958 127514 40010
rect 127566 39958 127618 40010
rect 158078 39958 158130 40010
rect 158182 39958 158234 40010
rect 158286 39958 158338 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 81278 39174 81330 39226
rect 81382 39174 81434 39226
rect 81486 39174 81538 39226
rect 111998 39174 112050 39226
rect 112102 39174 112154 39226
rect 112206 39174 112258 39226
rect 142718 39174 142770 39226
rect 142822 39174 142874 39226
rect 142926 39174 142978 39226
rect 173438 39174 173490 39226
rect 173542 39174 173594 39226
rect 173646 39174 173698 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 96638 38390 96690 38442
rect 96742 38390 96794 38442
rect 96846 38390 96898 38442
rect 127358 38390 127410 38442
rect 127462 38390 127514 38442
rect 127566 38390 127618 38442
rect 158078 38390 158130 38442
rect 158182 38390 158234 38442
rect 158286 38390 158338 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 81278 37606 81330 37658
rect 81382 37606 81434 37658
rect 81486 37606 81538 37658
rect 111998 37606 112050 37658
rect 112102 37606 112154 37658
rect 112206 37606 112258 37658
rect 142718 37606 142770 37658
rect 142822 37606 142874 37658
rect 142926 37606 142978 37658
rect 173438 37606 173490 37658
rect 173542 37606 173594 37658
rect 173646 37606 173698 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 96638 36822 96690 36874
rect 96742 36822 96794 36874
rect 96846 36822 96898 36874
rect 127358 36822 127410 36874
rect 127462 36822 127514 36874
rect 127566 36822 127618 36874
rect 158078 36822 158130 36874
rect 158182 36822 158234 36874
rect 158286 36822 158338 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 81278 36038 81330 36090
rect 81382 36038 81434 36090
rect 81486 36038 81538 36090
rect 111998 36038 112050 36090
rect 112102 36038 112154 36090
rect 112206 36038 112258 36090
rect 142718 36038 142770 36090
rect 142822 36038 142874 36090
rect 142926 36038 142978 36090
rect 173438 36038 173490 36090
rect 173542 36038 173594 36090
rect 173646 36038 173698 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 96638 35254 96690 35306
rect 96742 35254 96794 35306
rect 96846 35254 96898 35306
rect 127358 35254 127410 35306
rect 127462 35254 127514 35306
rect 127566 35254 127618 35306
rect 158078 35254 158130 35306
rect 158182 35254 158234 35306
rect 158286 35254 158338 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 81278 34470 81330 34522
rect 81382 34470 81434 34522
rect 81486 34470 81538 34522
rect 111998 34470 112050 34522
rect 112102 34470 112154 34522
rect 112206 34470 112258 34522
rect 142718 34470 142770 34522
rect 142822 34470 142874 34522
rect 142926 34470 142978 34522
rect 173438 34470 173490 34522
rect 173542 34470 173594 34522
rect 173646 34470 173698 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 96638 33686 96690 33738
rect 96742 33686 96794 33738
rect 96846 33686 96898 33738
rect 127358 33686 127410 33738
rect 127462 33686 127514 33738
rect 127566 33686 127618 33738
rect 158078 33686 158130 33738
rect 158182 33686 158234 33738
rect 158286 33686 158338 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 81278 32902 81330 32954
rect 81382 32902 81434 32954
rect 81486 32902 81538 32954
rect 111998 32902 112050 32954
rect 112102 32902 112154 32954
rect 112206 32902 112258 32954
rect 142718 32902 142770 32954
rect 142822 32902 142874 32954
rect 142926 32902 142978 32954
rect 173438 32902 173490 32954
rect 173542 32902 173594 32954
rect 173646 32902 173698 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 96638 32118 96690 32170
rect 96742 32118 96794 32170
rect 96846 32118 96898 32170
rect 127358 32118 127410 32170
rect 127462 32118 127514 32170
rect 127566 32118 127618 32170
rect 158078 32118 158130 32170
rect 158182 32118 158234 32170
rect 158286 32118 158338 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 81278 31334 81330 31386
rect 81382 31334 81434 31386
rect 81486 31334 81538 31386
rect 111998 31334 112050 31386
rect 112102 31334 112154 31386
rect 112206 31334 112258 31386
rect 142718 31334 142770 31386
rect 142822 31334 142874 31386
rect 142926 31334 142978 31386
rect 173438 31334 173490 31386
rect 173542 31334 173594 31386
rect 173646 31334 173698 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 96638 30550 96690 30602
rect 96742 30550 96794 30602
rect 96846 30550 96898 30602
rect 127358 30550 127410 30602
rect 127462 30550 127514 30602
rect 127566 30550 127618 30602
rect 158078 30550 158130 30602
rect 158182 30550 158234 30602
rect 158286 30550 158338 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 81278 29766 81330 29818
rect 81382 29766 81434 29818
rect 81486 29766 81538 29818
rect 111998 29766 112050 29818
rect 112102 29766 112154 29818
rect 112206 29766 112258 29818
rect 142718 29766 142770 29818
rect 142822 29766 142874 29818
rect 142926 29766 142978 29818
rect 173438 29766 173490 29818
rect 173542 29766 173594 29818
rect 173646 29766 173698 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 96638 28982 96690 29034
rect 96742 28982 96794 29034
rect 96846 28982 96898 29034
rect 127358 28982 127410 29034
rect 127462 28982 127514 29034
rect 127566 28982 127618 29034
rect 158078 28982 158130 29034
rect 158182 28982 158234 29034
rect 158286 28982 158338 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 81278 28198 81330 28250
rect 81382 28198 81434 28250
rect 81486 28198 81538 28250
rect 111998 28198 112050 28250
rect 112102 28198 112154 28250
rect 112206 28198 112258 28250
rect 142718 28198 142770 28250
rect 142822 28198 142874 28250
rect 142926 28198 142978 28250
rect 173438 28198 173490 28250
rect 173542 28198 173594 28250
rect 173646 28198 173698 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 96638 27414 96690 27466
rect 96742 27414 96794 27466
rect 96846 27414 96898 27466
rect 127358 27414 127410 27466
rect 127462 27414 127514 27466
rect 127566 27414 127618 27466
rect 158078 27414 158130 27466
rect 158182 27414 158234 27466
rect 158286 27414 158338 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 81278 26630 81330 26682
rect 81382 26630 81434 26682
rect 81486 26630 81538 26682
rect 111998 26630 112050 26682
rect 112102 26630 112154 26682
rect 112206 26630 112258 26682
rect 142718 26630 142770 26682
rect 142822 26630 142874 26682
rect 142926 26630 142978 26682
rect 173438 26630 173490 26682
rect 173542 26630 173594 26682
rect 173646 26630 173698 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 96638 25846 96690 25898
rect 96742 25846 96794 25898
rect 96846 25846 96898 25898
rect 127358 25846 127410 25898
rect 127462 25846 127514 25898
rect 127566 25846 127618 25898
rect 158078 25846 158130 25898
rect 158182 25846 158234 25898
rect 158286 25846 158338 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 81278 25062 81330 25114
rect 81382 25062 81434 25114
rect 81486 25062 81538 25114
rect 111998 25062 112050 25114
rect 112102 25062 112154 25114
rect 112206 25062 112258 25114
rect 142718 25062 142770 25114
rect 142822 25062 142874 25114
rect 142926 25062 142978 25114
rect 173438 25062 173490 25114
rect 173542 25062 173594 25114
rect 173646 25062 173698 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 96638 24278 96690 24330
rect 96742 24278 96794 24330
rect 96846 24278 96898 24330
rect 127358 24278 127410 24330
rect 127462 24278 127514 24330
rect 127566 24278 127618 24330
rect 158078 24278 158130 24330
rect 158182 24278 158234 24330
rect 158286 24278 158338 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 81278 23494 81330 23546
rect 81382 23494 81434 23546
rect 81486 23494 81538 23546
rect 111998 23494 112050 23546
rect 112102 23494 112154 23546
rect 112206 23494 112258 23546
rect 142718 23494 142770 23546
rect 142822 23494 142874 23546
rect 142926 23494 142978 23546
rect 173438 23494 173490 23546
rect 173542 23494 173594 23546
rect 173646 23494 173698 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 96638 22710 96690 22762
rect 96742 22710 96794 22762
rect 96846 22710 96898 22762
rect 127358 22710 127410 22762
rect 127462 22710 127514 22762
rect 127566 22710 127618 22762
rect 158078 22710 158130 22762
rect 158182 22710 158234 22762
rect 158286 22710 158338 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 81278 21926 81330 21978
rect 81382 21926 81434 21978
rect 81486 21926 81538 21978
rect 111998 21926 112050 21978
rect 112102 21926 112154 21978
rect 112206 21926 112258 21978
rect 142718 21926 142770 21978
rect 142822 21926 142874 21978
rect 142926 21926 142978 21978
rect 173438 21926 173490 21978
rect 173542 21926 173594 21978
rect 173646 21926 173698 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 96638 21142 96690 21194
rect 96742 21142 96794 21194
rect 96846 21142 96898 21194
rect 127358 21142 127410 21194
rect 127462 21142 127514 21194
rect 127566 21142 127618 21194
rect 158078 21142 158130 21194
rect 158182 21142 158234 21194
rect 158286 21142 158338 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 81278 20358 81330 20410
rect 81382 20358 81434 20410
rect 81486 20358 81538 20410
rect 111998 20358 112050 20410
rect 112102 20358 112154 20410
rect 112206 20358 112258 20410
rect 142718 20358 142770 20410
rect 142822 20358 142874 20410
rect 142926 20358 142978 20410
rect 173438 20358 173490 20410
rect 173542 20358 173594 20410
rect 173646 20358 173698 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 96638 19574 96690 19626
rect 96742 19574 96794 19626
rect 96846 19574 96898 19626
rect 127358 19574 127410 19626
rect 127462 19574 127514 19626
rect 127566 19574 127618 19626
rect 158078 19574 158130 19626
rect 158182 19574 158234 19626
rect 158286 19574 158338 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 81278 18790 81330 18842
rect 81382 18790 81434 18842
rect 81486 18790 81538 18842
rect 111998 18790 112050 18842
rect 112102 18790 112154 18842
rect 112206 18790 112258 18842
rect 142718 18790 142770 18842
rect 142822 18790 142874 18842
rect 142926 18790 142978 18842
rect 173438 18790 173490 18842
rect 173542 18790 173594 18842
rect 173646 18790 173698 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 96638 18006 96690 18058
rect 96742 18006 96794 18058
rect 96846 18006 96898 18058
rect 127358 18006 127410 18058
rect 127462 18006 127514 18058
rect 127566 18006 127618 18058
rect 158078 18006 158130 18058
rect 158182 18006 158234 18058
rect 158286 18006 158338 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 81278 17222 81330 17274
rect 81382 17222 81434 17274
rect 81486 17222 81538 17274
rect 111998 17222 112050 17274
rect 112102 17222 112154 17274
rect 112206 17222 112258 17274
rect 142718 17222 142770 17274
rect 142822 17222 142874 17274
rect 142926 17222 142978 17274
rect 173438 17222 173490 17274
rect 173542 17222 173594 17274
rect 173646 17222 173698 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 96638 16438 96690 16490
rect 96742 16438 96794 16490
rect 96846 16438 96898 16490
rect 127358 16438 127410 16490
rect 127462 16438 127514 16490
rect 127566 16438 127618 16490
rect 158078 16438 158130 16490
rect 158182 16438 158234 16490
rect 158286 16438 158338 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 81278 15654 81330 15706
rect 81382 15654 81434 15706
rect 81486 15654 81538 15706
rect 111998 15654 112050 15706
rect 112102 15654 112154 15706
rect 112206 15654 112258 15706
rect 142718 15654 142770 15706
rect 142822 15654 142874 15706
rect 142926 15654 142978 15706
rect 173438 15654 173490 15706
rect 173542 15654 173594 15706
rect 173646 15654 173698 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 96638 14870 96690 14922
rect 96742 14870 96794 14922
rect 96846 14870 96898 14922
rect 127358 14870 127410 14922
rect 127462 14870 127514 14922
rect 127566 14870 127618 14922
rect 158078 14870 158130 14922
rect 158182 14870 158234 14922
rect 158286 14870 158338 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 81278 14086 81330 14138
rect 81382 14086 81434 14138
rect 81486 14086 81538 14138
rect 111998 14086 112050 14138
rect 112102 14086 112154 14138
rect 112206 14086 112258 14138
rect 142718 14086 142770 14138
rect 142822 14086 142874 14138
rect 142926 14086 142978 14138
rect 173438 14086 173490 14138
rect 173542 14086 173594 14138
rect 173646 14086 173698 14138
rect 69134 13582 69186 13634
rect 69582 13582 69634 13634
rect 70030 13582 70082 13634
rect 70590 13582 70642 13634
rect 71038 13582 71090 13634
rect 72718 13582 72770 13634
rect 74958 13582 75010 13634
rect 75406 13582 75458 13634
rect 75854 13582 75906 13634
rect 77086 13582 77138 13634
rect 78206 13582 78258 13634
rect 79102 13582 79154 13634
rect 79774 13582 79826 13634
rect 80670 13582 80722 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 96638 13302 96690 13354
rect 96742 13302 96794 13354
rect 96846 13302 96898 13354
rect 127358 13302 127410 13354
rect 127462 13302 127514 13354
rect 127566 13302 127618 13354
rect 158078 13302 158130 13354
rect 158182 13302 158234 13354
rect 158286 13302 158338 13354
rect 75742 13134 75794 13186
rect 76414 13134 76466 13186
rect 79214 13134 79266 13186
rect 79550 13134 79602 13186
rect 79774 13134 79826 13186
rect 68238 13022 68290 13074
rect 69694 13022 69746 13074
rect 70142 13022 70194 13074
rect 71262 13022 71314 13074
rect 72270 13022 72322 13074
rect 73502 13022 73554 13074
rect 75742 13022 75794 13074
rect 83022 13022 83074 13074
rect 104078 13022 104130 13074
rect 76638 12910 76690 12962
rect 101166 12910 101218 12962
rect 79662 12798 79714 12850
rect 101950 12798 102002 12850
rect 67342 12686 67394 12738
rect 68686 12686 68738 12738
rect 70814 12686 70866 12738
rect 71710 12686 71762 12738
rect 72718 12686 72770 12738
rect 73166 12686 73218 12738
rect 74174 12686 74226 12738
rect 74734 12686 74786 12738
rect 75182 12686 75234 12738
rect 76190 12686 76242 12738
rect 77198 12686 77250 12738
rect 77758 12686 77810 12738
rect 78542 12686 78594 12738
rect 79102 12686 79154 12738
rect 79998 12686 80050 12738
rect 80894 12686 80946 12738
rect 81454 12686 81506 12738
rect 82686 12686 82738 12738
rect 100382 12686 100434 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 81278 12518 81330 12570
rect 81382 12518 81434 12570
rect 81486 12518 81538 12570
rect 111998 12518 112050 12570
rect 112102 12518 112154 12570
rect 112206 12518 112258 12570
rect 142718 12518 142770 12570
rect 142822 12518 142874 12570
rect 142926 12518 142978 12570
rect 173438 12518 173490 12570
rect 173542 12518 173594 12570
rect 173646 12518 173698 12570
rect 52782 12350 52834 12402
rect 57934 12350 57986 12402
rect 64206 12350 64258 12402
rect 70254 12350 70306 12402
rect 76078 12350 76130 12402
rect 76526 12350 76578 12402
rect 77086 12350 77138 12402
rect 77422 12350 77474 12402
rect 77982 12350 78034 12402
rect 79214 12350 79266 12402
rect 80558 12350 80610 12402
rect 81678 12350 81730 12402
rect 82574 12350 82626 12402
rect 85934 12350 85986 12402
rect 57374 12238 57426 12290
rect 59614 12238 59666 12290
rect 60846 12238 60898 12290
rect 61182 12238 61234 12290
rect 63758 12238 63810 12290
rect 73614 12238 73666 12290
rect 91086 12238 91138 12290
rect 91198 12126 91250 12178
rect 98814 12126 98866 12178
rect 105198 12126 105250 12178
rect 108670 12126 108722 12178
rect 55134 12014 55186 12066
rect 58382 12014 58434 12066
rect 59166 12014 59218 12066
rect 61966 12014 62018 12066
rect 64766 12014 64818 12066
rect 65662 12014 65714 12066
rect 66110 12014 66162 12066
rect 66894 12014 66946 12066
rect 67454 12014 67506 12066
rect 68126 12014 68178 12066
rect 68686 12014 68738 12066
rect 69134 12014 69186 12066
rect 69582 12014 69634 12066
rect 70590 12014 70642 12066
rect 71038 12014 71090 12066
rect 71934 12014 71986 12066
rect 72382 12014 72434 12066
rect 74174 12014 74226 12066
rect 74510 12014 74562 12066
rect 74958 12014 75010 12066
rect 75518 12014 75570 12066
rect 78542 12014 78594 12066
rect 79662 12014 79714 12066
rect 80110 12014 80162 12066
rect 81342 12014 81394 12066
rect 82238 12014 82290 12066
rect 83246 12014 83298 12066
rect 83694 12014 83746 12066
rect 84142 12014 84194 12066
rect 84814 12014 84866 12066
rect 90414 12014 90466 12066
rect 98142 12014 98194 12066
rect 99486 12014 99538 12066
rect 101614 12014 101666 12066
rect 104526 12014 104578 12066
rect 105982 12014 106034 12066
rect 108110 12014 108162 12066
rect 109454 12014 109506 12066
rect 111582 12014 111634 12066
rect 112142 12014 112194 12066
rect 57262 11902 57314 11954
rect 58382 11902 58434 11954
rect 60286 11902 60338 11954
rect 60622 11902 60674 11954
rect 68126 11902 68178 11954
rect 68574 11902 68626 11954
rect 91310 11902 91362 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 96638 11734 96690 11786
rect 96742 11734 96794 11786
rect 96846 11734 96898 11786
rect 127358 11734 127410 11786
rect 127462 11734 127514 11786
rect 127566 11734 127618 11786
rect 158078 11734 158130 11786
rect 158182 11734 158234 11786
rect 158286 11734 158338 11786
rect 57150 11566 57202 11618
rect 57934 11566 57986 11618
rect 99822 11566 99874 11618
rect 100606 11566 100658 11618
rect 47182 11454 47234 11506
rect 51998 11454 52050 11506
rect 54462 11454 54514 11506
rect 55022 11454 55074 11506
rect 57934 11454 57986 11506
rect 58382 11454 58434 11506
rect 59950 11454 60002 11506
rect 63758 11454 63810 11506
rect 67790 11454 67842 11506
rect 70142 11454 70194 11506
rect 77198 11454 77250 11506
rect 78094 11454 78146 11506
rect 79438 11454 79490 11506
rect 82798 11454 82850 11506
rect 85374 11454 85426 11506
rect 89518 11454 89570 11506
rect 91646 11454 91698 11506
rect 97246 11454 97298 11506
rect 99262 11454 99314 11506
rect 66558 11342 66610 11394
rect 69694 11342 69746 11394
rect 70702 11342 70754 11394
rect 72606 11342 72658 11394
rect 73390 11342 73442 11394
rect 78430 11342 78482 11394
rect 82238 11342 82290 11394
rect 88398 11342 88450 11394
rect 88958 11342 89010 11394
rect 92430 11342 92482 11394
rect 93774 11342 93826 11394
rect 94334 11330 94386 11382
rect 103406 11342 103458 11394
rect 106654 11342 106706 11394
rect 107438 11566 107490 11618
rect 107438 11454 107490 11506
rect 112030 11454 112082 11506
rect 115278 11454 115330 11506
rect 109118 11342 109170 11394
rect 51102 11230 51154 11282
rect 54014 11230 54066 11282
rect 65886 11230 65938 11282
rect 70814 11230 70866 11282
rect 71822 11230 71874 11282
rect 81566 11230 81618 11282
rect 83470 11230 83522 11282
rect 83694 11230 83746 11282
rect 87614 11230 87666 11282
rect 95118 11230 95170 11282
rect 99374 11230 99426 11282
rect 99934 11230 99986 11282
rect 104190 11230 104242 11282
rect 109902 11230 109954 11282
rect 39118 11118 39170 11170
rect 39566 11118 39618 11170
rect 46622 11118 46674 11170
rect 47630 11118 47682 11170
rect 48078 11118 48130 11170
rect 48750 11118 48802 11170
rect 51662 11118 51714 11170
rect 52782 11118 52834 11170
rect 53678 11118 53730 11170
rect 55582 11118 55634 11170
rect 56030 11118 56082 11170
rect 56366 11118 56418 11170
rect 56814 11118 56866 11170
rect 57486 11118 57538 11170
rect 58718 11118 58770 11170
rect 60286 11118 60338 11170
rect 61294 11118 61346 11170
rect 61854 11118 61906 11170
rect 62190 11118 62242 11170
rect 62638 11118 62690 11170
rect 63198 11118 63250 11170
rect 67118 11118 67170 11170
rect 68126 11118 68178 11170
rect 68574 11118 68626 11170
rect 69246 11118 69298 11170
rect 71038 11118 71090 11170
rect 71598 11118 71650 11170
rect 71710 11118 71762 11170
rect 75630 11118 75682 11170
rect 76190 11118 76242 11170
rect 78878 11118 78930 11170
rect 83582 11118 83634 11170
rect 84478 11118 84530 11170
rect 97694 11118 97746 11170
rect 98254 11118 98306 11170
rect 99150 11118 99202 11170
rect 100382 11118 100434 11170
rect 101166 11118 101218 11170
rect 101502 11118 101554 11170
rect 101950 11118 102002 11170
rect 102846 11118 102898 11170
rect 106430 11118 106482 11170
rect 107102 11118 107154 11170
rect 107886 11118 107938 11170
rect 108334 11118 108386 11170
rect 112702 11118 112754 11170
rect 113150 11118 113202 11170
rect 114718 11118 114770 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 81278 10950 81330 11002
rect 81382 10950 81434 11002
rect 81486 10950 81538 11002
rect 111998 10950 112050 11002
rect 112102 10950 112154 11002
rect 112206 10950 112258 11002
rect 142718 10950 142770 11002
rect 142822 10950 142874 11002
rect 142926 10950 142978 11002
rect 173438 10950 173490 11002
rect 173542 10950 173594 11002
rect 173646 10950 173698 11002
rect 39342 10782 39394 10834
rect 46398 10782 46450 10834
rect 48750 10782 48802 10834
rect 56030 10782 56082 10834
rect 63422 10782 63474 10834
rect 65550 10782 65602 10834
rect 74286 10782 74338 10834
rect 75742 10782 75794 10834
rect 76862 10782 76914 10834
rect 82126 10782 82178 10834
rect 86382 10782 86434 10834
rect 96462 10782 96514 10834
rect 100606 10782 100658 10834
rect 101054 10782 101106 10834
rect 101614 10782 101666 10834
rect 104302 10782 104354 10834
rect 105422 10782 105474 10834
rect 106430 10782 106482 10834
rect 108558 10782 108610 10834
rect 115054 10782 115106 10834
rect 115390 10782 115442 10834
rect 116734 10782 116786 10834
rect 37998 10670 38050 10722
rect 47630 10670 47682 10722
rect 51774 10670 51826 10722
rect 53230 10670 53282 10722
rect 57486 10670 57538 10722
rect 73950 10670 74002 10722
rect 74958 10670 75010 10722
rect 83470 10670 83522 10722
rect 103518 10670 103570 10722
rect 104190 10670 104242 10722
rect 105310 10670 105362 10722
rect 37774 10558 37826 10610
rect 42702 10558 42754 10610
rect 47854 10558 47906 10610
rect 52446 10558 52498 10610
rect 57822 10558 57874 10610
rect 61630 10558 61682 10610
rect 62302 10558 62354 10610
rect 68798 10558 68850 10610
rect 72494 10558 72546 10610
rect 73390 10558 73442 10610
rect 74846 10558 74898 10610
rect 75182 10558 75234 10610
rect 79774 10558 79826 10610
rect 81790 10558 81842 10610
rect 82686 10558 82738 10610
rect 86158 10558 86210 10610
rect 88174 10558 88226 10610
rect 92430 10558 92482 10610
rect 100158 10558 100210 10610
rect 109118 10558 109170 10610
rect 38782 10446 38834 10498
rect 39902 10446 39954 10498
rect 43374 10446 43426 10498
rect 45502 10446 45554 10498
rect 46062 10446 46114 10498
rect 47182 10446 47234 10498
rect 49870 10446 49922 10498
rect 50654 10446 50706 10498
rect 51214 10446 51266 10498
rect 55358 10446 55410 10498
rect 56478 10446 56530 10498
rect 58270 10446 58322 10498
rect 58830 10446 58882 10498
rect 59502 10446 59554 10498
rect 62862 10446 62914 10498
rect 63758 10446 63810 10498
rect 64206 10446 64258 10498
rect 64766 10446 64818 10498
rect 65998 10446 66050 10498
rect 68126 10446 68178 10498
rect 69694 10446 69746 10498
rect 71822 10446 71874 10498
rect 76190 10446 76242 10498
rect 79102 10446 79154 10498
rect 80446 10446 80498 10498
rect 81230 10446 81282 10498
rect 85598 10446 85650 10498
rect 87054 10446 87106 10498
rect 87614 10446 87666 10498
rect 88286 10446 88338 10498
rect 89518 10446 89570 10498
rect 91646 10446 91698 10498
rect 96014 10446 96066 10498
rect 97246 10446 97298 10498
rect 99374 10446 99426 10498
rect 101950 10446 102002 10498
rect 102398 10446 102450 10498
rect 102958 10446 103010 10498
rect 106094 10446 106146 10498
rect 106990 10446 107042 10498
rect 107326 10446 107378 10498
rect 108222 10446 108274 10498
rect 109902 10446 109954 10498
rect 112030 10446 112082 10498
rect 113150 10446 113202 10498
rect 113598 10446 113650 10498
rect 113934 10446 113986 10498
rect 114494 10446 114546 10498
rect 115950 10446 116002 10498
rect 117294 10446 117346 10498
rect 117742 10446 117794 10498
rect 118190 10446 118242 10498
rect 51662 10334 51714 10386
rect 58046 10334 58098 10386
rect 58270 10334 58322 10386
rect 58718 10334 58770 10386
rect 86494 10334 86546 10386
rect 88510 10334 88562 10386
rect 101278 10334 101330 10386
rect 101950 10334 102002 10386
rect 104414 10334 104466 10386
rect 105534 10334 105586 10386
rect 106542 10334 106594 10386
rect 107326 10334 107378 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 96638 10166 96690 10218
rect 96742 10166 96794 10218
rect 96846 10166 96898 10218
rect 127358 10166 127410 10218
rect 127462 10166 127514 10218
rect 127566 10166 127618 10218
rect 158078 10166 158130 10218
rect 158182 10166 158234 10218
rect 158286 10166 158338 10218
rect 51774 9998 51826 10050
rect 52670 9998 52722 10050
rect 54350 9998 54402 10050
rect 54686 9998 54738 10050
rect 61742 9998 61794 10050
rect 62078 9998 62130 10050
rect 83582 9998 83634 10050
rect 86942 9998 86994 10050
rect 87166 9998 87218 10050
rect 95454 9998 95506 10050
rect 104414 9998 104466 10050
rect 104638 9998 104690 10050
rect 106542 9998 106594 10050
rect 106990 9998 107042 10050
rect 114830 9998 114882 10050
rect 115502 9998 115554 10050
rect 118190 9998 118242 10050
rect 119086 9998 119138 10050
rect 33518 9886 33570 9938
rect 38334 9886 38386 9938
rect 40462 9886 40514 9938
rect 40910 9886 40962 9938
rect 43150 9886 43202 9938
rect 47406 9886 47458 9938
rect 49534 9886 49586 9938
rect 50878 9886 50930 9938
rect 53678 9886 53730 9938
rect 56926 9886 56978 9938
rect 59054 9886 59106 9938
rect 61742 9886 61794 9938
rect 62190 9886 62242 9938
rect 63422 9886 63474 9938
rect 63982 9886 64034 9938
rect 64766 9886 64818 9938
rect 73838 9886 73890 9938
rect 75294 9886 75346 9938
rect 76190 9886 76242 9938
rect 78654 9886 78706 9938
rect 84590 9886 84642 9938
rect 85822 9886 85874 9938
rect 86942 9886 86994 9938
rect 100270 9886 100322 9938
rect 103294 9886 103346 9938
rect 103630 9886 103682 9938
rect 104078 9886 104130 9938
rect 105198 9886 105250 9938
rect 106430 9886 106482 9938
rect 106990 9886 107042 9938
rect 108334 9886 108386 9938
rect 112142 9886 112194 9938
rect 113262 9886 113314 9938
rect 114158 9886 114210 9938
rect 116062 9886 116114 9938
rect 30718 9774 30770 9826
rect 37662 9774 37714 9826
rect 45614 9774 45666 9826
rect 46734 9774 46786 9826
rect 51438 9774 51490 9826
rect 52334 9774 52386 9826
rect 55470 9774 55522 9826
rect 56142 9774 56194 9826
rect 60174 9774 60226 9826
rect 68350 9774 68402 9826
rect 69358 9774 69410 9826
rect 77758 9774 77810 9826
rect 81006 9774 81058 9826
rect 81454 9774 81506 9826
rect 82238 9774 82290 9826
rect 88286 9774 88338 9826
rect 98142 9774 98194 9826
rect 98814 9774 98866 9826
rect 99150 9774 99202 9826
rect 102734 9774 102786 9826
rect 109230 9774 109282 9826
rect 117182 9774 117234 9826
rect 31390 9662 31442 9714
rect 36542 9662 36594 9714
rect 43710 9662 43762 9714
rect 44046 9662 44098 9714
rect 50430 9662 50482 9714
rect 55246 9662 55298 9714
rect 60510 9662 60562 9714
rect 67678 9662 67730 9714
rect 75182 9662 75234 9714
rect 76526 9662 76578 9714
rect 78766 9662 78818 9714
rect 79214 9662 79266 9714
rect 83918 9662 83970 9714
rect 87614 9662 87666 9714
rect 87726 9662 87778 9714
rect 89070 9662 89122 9714
rect 95790 9662 95842 9714
rect 96574 9662 96626 9714
rect 96910 9662 96962 9714
rect 97694 9662 97746 9714
rect 98366 9662 98418 9714
rect 101054 9662 101106 9714
rect 102398 9662 102450 9714
rect 110014 9662 110066 9714
rect 117070 9662 117122 9714
rect 117294 9662 117346 9714
rect 118526 9662 118578 9714
rect 119198 9662 119250 9714
rect 119422 9662 119474 9714
rect 33966 9550 34018 9602
rect 35198 9550 35250 9602
rect 36206 9550 36258 9602
rect 41470 9550 41522 9602
rect 42142 9550 42194 9602
rect 42590 9550 42642 9602
rect 44830 9550 44882 9602
rect 45838 9550 45890 9602
rect 50094 9550 50146 9602
rect 51662 9550 51714 9602
rect 52558 9550 52610 9602
rect 59614 9550 59666 9602
rect 62526 9550 62578 9602
rect 62974 9550 63026 9602
rect 64318 9550 64370 9602
rect 65438 9550 65490 9602
rect 75406 9550 75458 9602
rect 76302 9550 76354 9602
rect 77534 9550 77586 9602
rect 78542 9550 78594 9602
rect 79662 9550 79714 9602
rect 80110 9550 80162 9602
rect 80670 9550 80722 9602
rect 82574 9550 82626 9602
rect 83134 9550 83186 9602
rect 83694 9550 83746 9602
rect 85486 9550 85538 9602
rect 86494 9550 86546 9602
rect 87502 9550 87554 9602
rect 91310 9550 91362 9602
rect 95006 9550 95058 9602
rect 95566 9550 95618 9602
rect 97582 9550 97634 9602
rect 97918 9550 97970 9602
rect 99374 9550 99426 9602
rect 99486 9550 99538 9602
rect 99822 9550 99874 9602
rect 101502 9550 101554 9602
rect 104638 9550 104690 9602
rect 105534 9550 105586 9602
rect 105982 9550 106034 9602
rect 107438 9550 107490 9602
rect 107886 9550 107938 9602
rect 112814 9550 112866 9602
rect 113710 9550 113762 9602
rect 114718 9550 114770 9602
rect 115054 9550 115106 9602
rect 115502 9550 115554 9602
rect 118302 9550 118354 9602
rect 119870 9550 119922 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 81278 9382 81330 9434
rect 81382 9382 81434 9434
rect 81486 9382 81538 9434
rect 111998 9382 112050 9434
rect 112102 9382 112154 9434
rect 112206 9382 112258 9434
rect 142718 9382 142770 9434
rect 142822 9382 142874 9434
rect 142926 9382 142978 9434
rect 173438 9382 173490 9434
rect 173542 9382 173594 9434
rect 173646 9382 173698 9434
rect 31838 9214 31890 9266
rect 32846 9214 32898 9266
rect 35422 9214 35474 9266
rect 36990 9214 37042 9266
rect 41470 9214 41522 9266
rect 41918 9214 41970 9266
rect 42590 9214 42642 9266
rect 43038 9214 43090 9266
rect 43486 9214 43538 9266
rect 44606 9214 44658 9266
rect 46846 9214 46898 9266
rect 47518 9214 47570 9266
rect 55694 9214 55746 9266
rect 57934 9214 57986 9266
rect 65438 9214 65490 9266
rect 65774 9214 65826 9266
rect 66222 9214 66274 9266
rect 66894 9214 66946 9266
rect 67790 9214 67842 9266
rect 67902 9214 67954 9266
rect 68686 9214 68738 9266
rect 73726 9214 73778 9266
rect 74622 9214 74674 9266
rect 79662 9214 79714 9266
rect 80558 9214 80610 9266
rect 81566 9214 81618 9266
rect 88062 9214 88114 9266
rect 90190 9214 90242 9266
rect 94670 9214 94722 9266
rect 96238 9214 96290 9266
rect 99822 9214 99874 9266
rect 100494 9214 100546 9266
rect 100942 9214 100994 9266
rect 108558 9214 108610 9266
rect 113710 9214 113762 9266
rect 34638 9102 34690 9154
rect 45502 9102 45554 9154
rect 46510 9102 46562 9154
rect 48638 9102 48690 9154
rect 53566 9102 53618 9154
rect 55358 9102 55410 9154
rect 58606 9102 58658 9154
rect 58830 9102 58882 9154
rect 59614 9102 59666 9154
rect 71822 9102 71874 9154
rect 76078 9102 76130 9154
rect 89406 9102 89458 9154
rect 94782 9102 94834 9154
rect 95006 9102 95058 9154
rect 95118 9102 95170 9154
rect 96462 9102 96514 9154
rect 97358 9102 97410 9154
rect 99486 9102 99538 9154
rect 113038 9102 113090 9154
rect 32174 8990 32226 9042
rect 33742 8990 33794 9042
rect 34078 8990 34130 9042
rect 34526 8990 34578 9042
rect 37998 8990 38050 9042
rect 44942 8990 44994 9042
rect 45726 8990 45778 9042
rect 47854 8990 47906 9042
rect 48414 8990 48466 9042
rect 50318 8990 50370 9042
rect 56142 8990 56194 9042
rect 56702 8990 56754 9042
rect 60622 8990 60674 9042
rect 64430 8990 64482 9042
rect 72494 8990 72546 9042
rect 74510 8990 74562 9042
rect 75406 8990 75458 9042
rect 82126 8990 82178 9042
rect 83022 8990 83074 9042
rect 86494 8990 86546 9042
rect 89294 8990 89346 9042
rect 89630 8990 89682 9042
rect 93214 8990 93266 9042
rect 95902 8990 95954 9042
rect 98366 8990 98418 9042
rect 98814 8990 98866 9042
rect 99710 8990 99762 9042
rect 100158 8990 100210 9042
rect 104302 8990 104354 9042
rect 105198 8990 105250 9042
rect 109118 8990 109170 9042
rect 35870 8878 35922 8930
rect 36318 8878 36370 8930
rect 37438 8878 37490 8930
rect 38670 8878 38722 8930
rect 40798 8878 40850 8930
rect 44046 8878 44098 8930
rect 58270 8878 58322 8930
rect 61294 8878 61346 8930
rect 63422 8878 63474 8930
rect 64206 8878 64258 8930
rect 66782 8878 66834 8930
rect 68574 8878 68626 8930
rect 69694 8878 69746 8930
rect 73614 8878 73666 8930
rect 78206 8878 78258 8930
rect 78766 8878 78818 8930
rect 80110 8878 80162 8930
rect 83582 8878 83634 8930
rect 85710 8878 85762 8930
rect 86942 8878 86994 8930
rect 87614 8878 87666 8930
rect 88510 8878 88562 8930
rect 92430 8878 92482 8930
rect 94222 8878 94274 8930
rect 98926 8878 98978 8930
rect 101502 8878 101554 8930
rect 103630 8878 103682 8930
rect 105982 8878 106034 8930
rect 108110 8878 108162 8930
rect 109902 8878 109954 8930
rect 112030 8878 112082 8930
rect 113486 8878 113538 8930
rect 35758 8766 35810 8818
rect 36318 8766 36370 8818
rect 64094 8766 64146 8818
rect 67118 8766 67170 8818
rect 68014 8766 68066 8818
rect 68910 8766 68962 8818
rect 73950 8766 74002 8818
rect 74622 8766 74674 8818
rect 78878 8766 78930 8818
rect 82126 8766 82178 8818
rect 82462 8766 82514 8818
rect 95230 8766 95282 8818
rect 96574 8766 96626 8818
rect 114382 9214 114434 9266
rect 114830 9214 114882 9266
rect 116622 9214 116674 9266
rect 118638 9214 118690 9266
rect 120990 9214 121042 9266
rect 121886 9214 121938 9266
rect 115390 9102 115442 9154
rect 115726 9102 115778 9154
rect 116286 9102 116338 9154
rect 117182 9102 117234 9154
rect 117518 9102 117570 9154
rect 114046 8990 114098 9042
rect 118414 8990 118466 9042
rect 121550 8990 121602 9042
rect 119198 8878 119250 8930
rect 119646 8878 119698 8930
rect 120094 8878 120146 8930
rect 97246 8766 97298 8818
rect 113822 8766 113874 8818
rect 118750 8766 118802 8818
rect 119534 8766 119586 8818
rect 120094 8766 120146 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 96638 8598 96690 8650
rect 96742 8598 96794 8650
rect 96846 8598 96898 8650
rect 127358 8598 127410 8650
rect 127462 8598 127514 8650
rect 127566 8598 127618 8650
rect 158078 8598 158130 8650
rect 158182 8598 158234 8650
rect 158286 8598 158338 8650
rect 38222 8430 38274 8482
rect 42478 8430 42530 8482
rect 43150 8430 43202 8482
rect 59726 8430 59778 8482
rect 60062 8430 60114 8482
rect 94782 8430 94834 8482
rect 98814 8430 98866 8482
rect 33630 8318 33682 8370
rect 37886 8318 37938 8370
rect 40126 8318 40178 8370
rect 43038 8318 43090 8370
rect 43934 8318 43986 8370
rect 48190 8318 48242 8370
rect 50318 8318 50370 8370
rect 55246 8318 55298 8370
rect 60174 8318 60226 8370
rect 68238 8318 68290 8370
rect 68574 8318 68626 8370
rect 73502 8318 73554 8370
rect 78542 8318 78594 8370
rect 82462 8318 82514 8370
rect 83694 8318 83746 8370
rect 85710 8318 85762 8370
rect 86270 8318 86322 8370
rect 90302 8318 90354 8370
rect 91870 8318 91922 8370
rect 92430 8318 92482 8370
rect 93774 8318 93826 8370
rect 94222 8318 94274 8370
rect 100382 8430 100434 8482
rect 95342 8318 95394 8370
rect 100046 8318 100098 8370
rect 100158 8318 100210 8370
rect 101838 8318 101890 8370
rect 105198 8318 105250 8370
rect 113262 8318 113314 8370
rect 117518 8318 117570 8370
rect 123454 8318 123506 8370
rect 138798 8318 138850 8370
rect 30718 8206 30770 8258
rect 35086 8206 35138 8258
rect 38894 8206 38946 8258
rect 45502 8206 45554 8258
rect 50990 8206 51042 8258
rect 51886 8206 51938 8258
rect 52110 8206 52162 8258
rect 52446 8206 52498 8258
rect 53342 8206 53394 8258
rect 54014 8206 54066 8258
rect 54798 8206 54850 8258
rect 59278 8206 59330 8258
rect 61406 8206 61458 8258
rect 67342 8206 67394 8258
rect 69358 8206 69410 8258
rect 75406 8206 75458 8258
rect 77422 8206 77474 8258
rect 78990 8206 79042 8258
rect 80670 8206 80722 8258
rect 80894 8206 80946 8258
rect 81118 8206 81170 8258
rect 82574 8206 82626 8258
rect 84254 8206 84306 8258
rect 84590 8206 84642 8258
rect 85486 8206 85538 8258
rect 87278 8206 87330 8258
rect 87502 8206 87554 8258
rect 90190 8206 90242 8258
rect 91646 8206 91698 8258
rect 94894 8206 94946 8258
rect 95566 8206 95618 8258
rect 96350 8206 96402 8258
rect 97806 8206 97858 8258
rect 98590 8206 98642 8258
rect 99150 8206 99202 8258
rect 99486 8206 99538 8258
rect 101390 8206 101442 8258
rect 102846 8206 102898 8258
rect 103742 8206 103794 8258
rect 104414 8206 104466 8258
rect 108334 8206 108386 8258
rect 109342 8206 109394 8258
rect 114942 8206 114994 8258
rect 116062 8206 116114 8258
rect 116958 8206 117010 8258
rect 119646 8206 119698 8258
rect 119758 8206 119810 8258
rect 120654 8206 120706 8258
rect 19630 8094 19682 8146
rect 27134 8094 27186 8146
rect 31502 8094 31554 8146
rect 34302 8094 34354 8146
rect 34750 8094 34802 8146
rect 36430 8094 36482 8146
rect 39006 8094 39058 8146
rect 40350 8094 40402 8146
rect 40798 8094 40850 8146
rect 46398 8094 46450 8146
rect 46734 8094 46786 8146
rect 47294 8094 47346 8146
rect 53790 8094 53842 8146
rect 56254 8094 56306 8146
rect 57486 8094 57538 8146
rect 57822 8094 57874 8146
rect 66446 8094 66498 8146
rect 75518 8094 75570 8146
rect 76190 8094 76242 8146
rect 76526 8094 76578 8146
rect 78206 8094 78258 8146
rect 78430 8094 78482 8146
rect 79326 8094 79378 8146
rect 79886 8094 79938 8146
rect 81342 8094 81394 8146
rect 83246 8094 83298 8146
rect 85262 8094 85314 8146
rect 85822 8094 85874 8146
rect 86718 8094 86770 8146
rect 87838 8094 87890 8146
rect 88734 8094 88786 8146
rect 91086 8094 91138 8146
rect 91982 8094 92034 8146
rect 96686 8094 96738 8146
rect 98030 8094 98082 8146
rect 98142 8094 98194 8146
rect 99710 8094 99762 8146
rect 99822 8094 99874 8146
rect 101614 8094 101666 8146
rect 101950 8094 102002 8146
rect 103966 8094 104018 8146
rect 105310 8094 105362 8146
rect 107214 8094 107266 8146
rect 110014 8094 110066 8146
rect 113710 8094 113762 8146
rect 119534 8094 119586 8146
rect 19294 7982 19346 8034
rect 26798 7982 26850 8034
rect 27806 7982 27858 8034
rect 28814 7982 28866 8034
rect 29598 7982 29650 8034
rect 35422 7982 35474 8034
rect 36878 7982 36930 8034
rect 39790 7982 39842 8034
rect 41806 7982 41858 8034
rect 42254 7982 42306 8034
rect 42590 7982 42642 8034
rect 43710 7982 43762 8034
rect 43822 7982 43874 8034
rect 44830 7982 44882 8034
rect 45838 7982 45890 8034
rect 47630 7982 47682 8034
rect 52334 7982 52386 8034
rect 53566 7982 53618 8034
rect 55918 7982 55970 8034
rect 57038 7982 57090 8034
rect 58382 7982 58434 8034
rect 58942 7982 58994 8034
rect 59726 7982 59778 8034
rect 60734 7982 60786 8034
rect 67678 7982 67730 8034
rect 75742 7982 75794 8034
rect 77646 7982 77698 8034
rect 79214 7982 79266 8034
rect 80222 7982 80274 8034
rect 84366 7982 84418 8034
rect 88398 7982 88450 8034
rect 89406 7982 89458 8034
rect 93102 7982 93154 8034
rect 95678 7982 95730 8034
rect 96238 7982 96290 8034
rect 96462 7982 96514 8034
rect 97246 7982 97298 8034
rect 102398 7982 102450 8034
rect 105086 7982 105138 8034
rect 105758 7982 105810 8034
rect 106206 7982 106258 8034
rect 106654 7982 106706 8034
rect 107998 7982 108050 8034
rect 112254 7982 112306 8034
rect 112814 7982 112866 8034
rect 114158 7982 114210 8034
rect 115166 7982 115218 8034
rect 115726 7982 115778 8034
rect 117854 7982 117906 8034
rect 118302 7982 118354 8034
rect 118862 7982 118914 8034
rect 120206 7982 120258 8034
rect 121102 7982 121154 8034
rect 121550 7982 121602 8034
rect 121998 7982 122050 8034
rect 122558 7982 122610 8034
rect 123006 7982 123058 8034
rect 123790 7982 123842 8034
rect 124350 7982 124402 8034
rect 128830 7982 128882 8034
rect 130622 7982 130674 8034
rect 131070 7982 131122 8034
rect 131406 7982 131458 8034
rect 131966 7982 132018 8034
rect 132974 7982 133026 8034
rect 133646 7982 133698 8034
rect 135102 7982 135154 8034
rect 135438 7982 135490 8034
rect 136670 7982 136722 8034
rect 137566 7982 137618 8034
rect 139694 7982 139746 8034
rect 140142 7982 140194 8034
rect 140926 7982 140978 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 81278 7814 81330 7866
rect 81382 7814 81434 7866
rect 81486 7814 81538 7866
rect 111998 7814 112050 7866
rect 112102 7814 112154 7866
rect 112206 7814 112258 7866
rect 142718 7814 142770 7866
rect 142822 7814 142874 7866
rect 142926 7814 142978 7866
rect 173438 7814 173490 7866
rect 173542 7814 173594 7866
rect 173646 7814 173698 7866
rect 31950 7646 32002 7698
rect 37886 7646 37938 7698
rect 39230 7646 39282 7698
rect 47294 7646 47346 7698
rect 55694 7646 55746 7698
rect 61742 7646 61794 7698
rect 62414 7646 62466 7698
rect 73390 7646 73442 7698
rect 75406 7646 75458 7698
rect 80110 7646 80162 7698
rect 81678 7646 81730 7698
rect 90862 7646 90914 7698
rect 91758 7646 91810 7698
rect 93102 7646 93154 7698
rect 93550 7646 93602 7698
rect 93998 7646 94050 7698
rect 94446 7646 94498 7698
rect 94894 7646 94946 7698
rect 97806 7646 97858 7698
rect 98366 7646 98418 7698
rect 99710 7646 99762 7698
rect 100046 7646 100098 7698
rect 100942 7646 100994 7698
rect 101502 7646 101554 7698
rect 102398 7646 102450 7698
rect 103406 7646 103458 7698
rect 103518 7646 103570 7698
rect 104302 7646 104354 7698
rect 105534 7646 105586 7698
rect 106878 7646 106930 7698
rect 107438 7646 107490 7698
rect 109566 7646 109618 7698
rect 109902 7646 109954 7698
rect 112366 7646 112418 7698
rect 114382 7646 114434 7698
rect 114830 7646 114882 7698
rect 115838 7646 115890 7698
rect 120990 7646 121042 7698
rect 123230 7646 123282 7698
rect 124238 7646 124290 7698
rect 129950 7646 130002 7698
rect 130846 7646 130898 7698
rect 131518 7646 131570 7698
rect 132414 7646 132466 7698
rect 134430 7646 134482 7698
rect 137790 7646 137842 7698
rect 138798 7646 138850 7698
rect 18958 7534 19010 7586
rect 26462 7534 26514 7586
rect 32286 7534 32338 7586
rect 39566 7534 39618 7586
rect 42814 7534 42866 7586
rect 44158 7534 44210 7586
rect 51102 7534 51154 7586
rect 56030 7534 56082 7586
rect 56254 7534 56306 7586
rect 62862 7534 62914 7586
rect 69022 7534 69074 7586
rect 73726 7534 73778 7586
rect 74286 7534 74338 7586
rect 76526 7534 76578 7586
rect 78990 7534 79042 7586
rect 81566 7534 81618 7586
rect 83918 7534 83970 7586
rect 85038 7534 85090 7586
rect 95006 7534 95058 7586
rect 95230 7534 95282 7586
rect 95678 7534 95730 7586
rect 97358 7534 97410 7586
rect 101838 7534 101890 7586
rect 104190 7534 104242 7586
rect 107998 7534 108050 7586
rect 108110 7534 108162 7586
rect 113150 7534 113202 7586
rect 115950 7534 116002 7586
rect 117630 7534 117682 7586
rect 118190 7534 118242 7586
rect 118414 7534 118466 7586
rect 121438 7534 121490 7586
rect 18286 7422 18338 7474
rect 25678 7422 25730 7474
rect 33518 7422 33570 7474
rect 34190 7422 34242 7474
rect 36094 7422 36146 7474
rect 37550 7422 37602 7474
rect 42478 7422 42530 7474
rect 43374 7422 43426 7474
rect 46958 7422 47010 7474
rect 47854 7422 47906 7474
rect 53902 7422 53954 7474
rect 55358 7422 55410 7474
rect 56366 7422 56418 7474
rect 56702 7422 56754 7474
rect 57822 7422 57874 7474
rect 62302 7422 62354 7474
rect 62526 7422 62578 7474
rect 63422 7422 63474 7474
rect 63646 7422 63698 7474
rect 63870 7422 63922 7474
rect 66894 7422 66946 7474
rect 71598 7422 71650 7474
rect 74510 7422 74562 7474
rect 75294 7422 75346 7474
rect 76414 7422 76466 7474
rect 78542 7422 78594 7474
rect 82350 7422 82402 7474
rect 84814 7422 84866 7474
rect 86830 7422 86882 7474
rect 89518 7422 89570 7474
rect 89854 7422 89906 7474
rect 95454 7422 95506 7474
rect 100494 7422 100546 7474
rect 102734 7422 102786 7474
rect 106430 7422 106482 7474
rect 107774 7422 107826 7474
rect 110798 7422 110850 7474
rect 112030 7422 112082 7474
rect 113374 7422 113426 7474
rect 115390 7422 115442 7474
rect 115614 7422 115666 7474
rect 117294 7422 117346 7474
rect 118750 7422 118802 7474
rect 119646 7422 119698 7474
rect 130398 7422 130450 7474
rect 131966 7422 132018 7474
rect 14926 7310 14978 7362
rect 16382 7310 16434 7362
rect 21086 7310 21138 7362
rect 21534 7310 21586 7362
rect 21982 7310 22034 7362
rect 22430 7310 22482 7362
rect 22878 7310 22930 7362
rect 23438 7310 23490 7362
rect 23886 7310 23938 7362
rect 24222 7310 24274 7362
rect 28590 7310 28642 7362
rect 29038 7310 29090 7362
rect 29598 7310 29650 7362
rect 30046 7310 30098 7362
rect 30606 7310 30658 7362
rect 30942 7310 30994 7362
rect 31502 7310 31554 7362
rect 32846 7310 32898 7362
rect 34638 7310 34690 7362
rect 35310 7310 35362 7362
rect 36654 7310 36706 7362
rect 36990 7310 37042 7362
rect 38782 7310 38834 7362
rect 40462 7310 40514 7362
rect 40910 7310 40962 7362
rect 41582 7310 41634 7362
rect 41918 7310 41970 7362
rect 46286 7310 46338 7362
rect 48414 7310 48466 7362
rect 58606 7310 58658 7362
rect 60734 7310 60786 7362
rect 61406 7310 61458 7362
rect 63534 7310 63586 7362
rect 64654 7310 64706 7362
rect 71710 7310 71762 7362
rect 83134 7310 83186 7362
rect 86494 7310 86546 7362
rect 87278 7310 87330 7362
rect 87726 7310 87778 7362
rect 88510 7310 88562 7362
rect 90414 7310 90466 7362
rect 92094 7310 92146 7362
rect 92766 7310 92818 7362
rect 96126 7310 96178 7362
rect 97246 7310 97298 7362
rect 98702 7310 98754 7362
rect 99150 7310 99202 7362
rect 105086 7310 105138 7362
rect 105982 7310 106034 7362
rect 108558 7310 108610 7362
rect 109006 7310 109058 7362
rect 110350 7310 110402 7362
rect 111246 7310 111298 7362
rect 113934 7310 113986 7362
rect 116398 7310 116450 7362
rect 118638 7310 118690 7362
rect 119422 7310 119474 7362
rect 120318 7310 120370 7362
rect 121998 7310 122050 7362
rect 122446 7310 122498 7362
rect 122894 7310 122946 7362
rect 123790 7310 123842 7362
rect 124686 7310 124738 7362
rect 125022 7310 125074 7362
rect 125470 7310 125522 7362
rect 126142 7310 126194 7362
rect 126478 7310 126530 7362
rect 127934 7310 127986 7362
rect 128382 7310 128434 7362
rect 128942 7310 128994 7362
rect 129502 7310 129554 7362
rect 132750 7310 132802 7362
rect 133198 7310 133250 7362
rect 134094 7310 134146 7362
rect 135214 7310 135266 7362
rect 135662 7310 135714 7362
rect 136110 7310 136162 7362
rect 136894 7310 136946 7362
rect 137342 7310 137394 7362
rect 138238 7310 138290 7362
rect 139134 7310 139186 7362
rect 140030 7310 140082 7362
rect 140478 7310 140530 7362
rect 140926 7310 140978 7362
rect 141598 7310 141650 7362
rect 141934 7310 141986 7362
rect 142718 7310 142770 7362
rect 143054 7310 143106 7362
rect 143614 7310 143666 7362
rect 144846 7310 144898 7362
rect 145406 7310 145458 7362
rect 35758 7198 35810 7250
rect 36094 7198 36146 7250
rect 56702 7198 56754 7250
rect 72382 7198 72434 7250
rect 75406 7198 75458 7250
rect 81678 7198 81730 7250
rect 103294 7198 103346 7250
rect 109342 7198 109394 7250
rect 110014 7198 110066 7250
rect 124462 7198 124514 7250
rect 124686 7198 124738 7250
rect 132862 7198 132914 7250
rect 133198 7198 133250 7250
rect 136782 7198 136834 7250
rect 137790 7198 137842 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 96638 7030 96690 7082
rect 96742 7030 96794 7082
rect 96846 7030 96898 7082
rect 127358 7030 127410 7082
rect 127462 7030 127514 7082
rect 127566 7030 127618 7082
rect 158078 7030 158130 7082
rect 158182 7030 158234 7082
rect 158286 7030 158338 7082
rect 19630 6862 19682 6914
rect 19966 6862 20018 6914
rect 27470 6862 27522 6914
rect 45950 6862 46002 6914
rect 50430 6862 50482 6914
rect 77758 6862 77810 6914
rect 83134 6862 83186 6914
rect 83470 6862 83522 6914
rect 87502 6862 87554 6914
rect 87726 6862 87778 6914
rect 91198 6862 91250 6914
rect 91758 6862 91810 6914
rect 135774 6862 135826 6914
rect 141598 6862 141650 6914
rect 142158 6862 142210 6914
rect 143054 6862 143106 6914
rect 143838 6862 143890 6914
rect 27806 6750 27858 6802
rect 32062 6750 32114 6802
rect 56366 6750 56418 6802
rect 62974 6750 63026 6802
rect 65102 6750 65154 6802
rect 73838 6750 73890 6802
rect 76526 6750 76578 6802
rect 77534 6750 77586 6802
rect 80670 6750 80722 6802
rect 85822 6750 85874 6802
rect 87726 6750 87778 6802
rect 89742 6750 89794 6802
rect 95118 6750 95170 6802
rect 96686 6750 96738 6802
rect 97358 6750 97410 6802
rect 101502 6750 101554 6802
rect 102734 6750 102786 6802
rect 105870 6750 105922 6802
rect 109342 6750 109394 6802
rect 114382 6750 114434 6802
rect 115502 6750 115554 6802
rect 119086 6750 119138 6802
rect 120206 6750 120258 6802
rect 122894 6750 122946 6802
rect 20638 6638 20690 6690
rect 24110 6638 24162 6690
rect 25902 6638 25954 6690
rect 34862 6638 34914 6690
rect 35982 6638 36034 6690
rect 36430 6638 36482 6690
rect 37438 6638 37490 6690
rect 37774 6638 37826 6690
rect 38894 6638 38946 6690
rect 42366 6638 42418 6690
rect 42926 6638 42978 6690
rect 43374 6638 43426 6690
rect 44606 6638 44658 6690
rect 45614 6638 45666 6690
rect 46734 6638 46786 6690
rect 49758 6638 49810 6690
rect 50766 6638 50818 6690
rect 51438 6638 51490 6690
rect 53454 6638 53506 6690
rect 54238 6638 54290 6690
rect 57150 6638 57202 6690
rect 62190 6638 62242 6690
rect 65886 6638 65938 6690
rect 66110 6638 66162 6690
rect 66334 6638 66386 6690
rect 66558 6638 66610 6690
rect 68574 6638 68626 6690
rect 69358 6638 69410 6690
rect 77310 6638 77362 6690
rect 79662 6638 79714 6690
rect 80782 6638 80834 6690
rect 82126 6638 82178 6690
rect 82910 6638 82962 6690
rect 85262 6638 85314 6690
rect 87278 6638 87330 6690
rect 89294 6638 89346 6690
rect 91534 6638 91586 6690
rect 91982 6638 92034 6690
rect 92318 6638 92370 6690
rect 93102 6638 93154 6690
rect 93774 6638 93826 6690
rect 95678 6638 95730 6690
rect 95902 6638 95954 6690
rect 96238 6638 96290 6690
rect 97470 6638 97522 6690
rect 97694 6638 97746 6690
rect 99486 6638 99538 6690
rect 99934 6638 99986 6690
rect 101054 6638 101106 6690
rect 102622 6638 102674 6690
rect 103966 6638 104018 6690
rect 104190 6638 104242 6690
rect 105086 6638 105138 6690
rect 106766 6638 106818 6690
rect 110238 6638 110290 6690
rect 111134 6638 111186 6690
rect 112142 6638 112194 6690
rect 113934 6638 113986 6690
rect 117406 6638 117458 6690
rect 119310 6638 119362 6690
rect 120430 6638 120482 6690
rect 122446 6638 122498 6690
rect 123902 6638 123954 6690
rect 126926 6638 126978 6690
rect 128046 6638 128098 6690
rect 128606 6638 128658 6690
rect 128942 6638 128994 6690
rect 130062 6638 130114 6690
rect 130622 6638 130674 6690
rect 130958 6638 131010 6690
rect 132302 6638 132354 6690
rect 135886 6638 135938 6690
rect 141262 6638 141314 6690
rect 143950 6638 144002 6690
rect 14590 6526 14642 6578
rect 18734 6526 18786 6578
rect 20750 6526 20802 6578
rect 21534 6526 21586 6578
rect 22654 6526 22706 6578
rect 24334 6526 24386 6578
rect 28142 6526 28194 6578
rect 28590 6526 28642 6578
rect 29598 6526 29650 6578
rect 29934 6526 29986 6578
rect 30494 6526 30546 6578
rect 34190 6526 34242 6578
rect 35758 6526 35810 6578
rect 36206 6526 36258 6578
rect 38110 6526 38162 6578
rect 39678 6526 39730 6578
rect 40014 6526 40066 6578
rect 40574 6526 40626 6578
rect 40910 6526 40962 6578
rect 41806 6526 41858 6578
rect 42590 6526 42642 6578
rect 42814 6526 42866 6578
rect 44382 6526 44434 6578
rect 46510 6526 46562 6578
rect 47742 6526 47794 6578
rect 48078 6526 48130 6578
rect 48638 6526 48690 6578
rect 48974 6526 49026 6578
rect 49646 6526 49698 6578
rect 52334 6526 52386 6578
rect 57710 6526 57762 6578
rect 58046 6526 58098 6578
rect 59390 6526 59442 6578
rect 60622 6526 60674 6578
rect 67678 6526 67730 6578
rect 68126 6526 68178 6578
rect 75518 6526 75570 6578
rect 78430 6526 78482 6578
rect 78766 6526 78818 6578
rect 79774 6526 79826 6578
rect 81454 6526 81506 6578
rect 82238 6526 82290 6578
rect 84478 6526 84530 6578
rect 85822 6526 85874 6578
rect 86830 6526 86882 6578
rect 97246 6526 97298 6578
rect 98590 6526 98642 6578
rect 99038 6526 99090 6578
rect 103070 6526 103122 6578
rect 104526 6526 104578 6578
rect 105646 6526 105698 6578
rect 106654 6526 106706 6578
rect 109118 6526 109170 6578
rect 113038 6526 113090 6578
rect 115726 6526 115778 6578
rect 115950 6526 116002 6578
rect 116062 6526 116114 6578
rect 117854 6526 117906 6578
rect 121102 6526 121154 6578
rect 129726 6526 129778 6578
rect 136670 6526 136722 6578
rect 139134 6526 139186 6578
rect 14142 6414 14194 6466
rect 14926 6414 14978 6466
rect 15486 6414 15538 6466
rect 15822 6414 15874 6466
rect 16382 6414 16434 6466
rect 16942 6414 16994 6466
rect 17390 6414 17442 6466
rect 17726 6414 17778 6466
rect 18174 6414 18226 6466
rect 18846 6414 18898 6466
rect 19070 6414 19122 6466
rect 22206 6414 22258 6466
rect 23214 6414 23266 6466
rect 24782 6414 24834 6466
rect 25342 6414 25394 6466
rect 26126 6414 26178 6466
rect 26910 6414 26962 6466
rect 31054 6414 31106 6466
rect 31614 6414 31666 6466
rect 36878 6414 36930 6466
rect 37774 6414 37826 6466
rect 39118 6414 39170 6466
rect 41470 6414 41522 6466
rect 43822 6414 43874 6466
rect 58830 6414 58882 6466
rect 59726 6414 59778 6466
rect 60398 6414 60450 6466
rect 60510 6414 60562 6466
rect 61742 6414 61794 6466
rect 67006 6414 67058 6466
rect 67902 6414 67954 6466
rect 68238 6414 68290 6466
rect 75182 6414 75234 6466
rect 76414 6414 76466 6466
rect 77422 6414 77474 6466
rect 79998 6414 80050 6466
rect 82462 6414 82514 6466
rect 84142 6414 84194 6466
rect 85486 6414 85538 6466
rect 85710 6414 85762 6466
rect 86494 6414 86546 6466
rect 88398 6414 88450 6466
rect 90078 6414 90130 6466
rect 90526 6414 90578 6466
rect 90974 6414 91026 6466
rect 94446 6414 94498 6466
rect 95902 6414 95954 6466
rect 98254 6414 98306 6466
rect 100382 6414 100434 6466
rect 109342 6414 109394 6466
rect 110574 6414 110626 6466
rect 111246 6414 111298 6466
rect 111694 6414 111746 6466
rect 112590 6414 112642 6466
rect 113486 6414 113538 6466
rect 114830 6414 114882 6466
rect 116286 6414 116338 6466
rect 117070 6414 117122 6466
rect 118750 6414 118802 6466
rect 121550 6414 121602 6466
rect 121998 6414 122050 6466
rect 123454 6414 123506 6466
rect 124238 6414 124290 6466
rect 124910 6414 124962 6466
rect 125358 6414 125410 6466
rect 125806 6414 125858 6466
rect 126478 6414 126530 6466
rect 127374 6414 127426 6466
rect 129838 6414 129890 6466
rect 130734 6414 130786 6466
rect 131630 6414 131682 6466
rect 133310 6414 133362 6466
rect 133870 6414 133922 6466
rect 134318 6414 134370 6466
rect 134990 6414 135042 6466
rect 135998 6414 136050 6466
rect 137230 6414 137282 6466
rect 137678 6414 137730 6466
rect 138126 6414 138178 6466
rect 138686 6414 138738 6466
rect 139582 6414 139634 6466
rect 139918 6414 139970 6466
rect 140926 6414 140978 6466
rect 141710 6414 141762 6466
rect 142270 6414 142322 6466
rect 142606 6414 142658 6466
rect 143054 6414 143106 6466
rect 143502 6414 143554 6466
rect 144510 6414 144562 6466
rect 145070 6414 145122 6466
rect 145742 6414 145794 6466
rect 146302 6414 146354 6466
rect 146638 6414 146690 6466
rect 147086 6414 147138 6466
rect 147646 6414 147698 6466
rect 148766 6414 148818 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 81278 6246 81330 6298
rect 81382 6246 81434 6298
rect 81486 6246 81538 6298
rect 111998 6246 112050 6298
rect 112102 6246 112154 6298
rect 112206 6246 112258 6298
rect 142718 6246 142770 6298
rect 142822 6246 142874 6298
rect 142926 6246 142978 6298
rect 173438 6246 173490 6298
rect 173542 6246 173594 6298
rect 173646 6246 173698 6298
rect 15262 6078 15314 6130
rect 16046 6078 16098 6130
rect 16718 6078 16770 6130
rect 16942 6078 16994 6130
rect 22766 6078 22818 6130
rect 23550 6078 23602 6130
rect 24446 6078 24498 6130
rect 24894 6078 24946 6130
rect 29150 6078 29202 6130
rect 32846 6078 32898 6130
rect 34974 6078 35026 6130
rect 39342 6078 39394 6130
rect 41918 6078 41970 6130
rect 46062 6078 46114 6130
rect 46846 6078 46898 6130
rect 47742 6078 47794 6130
rect 56590 6078 56642 6130
rect 59390 6078 59442 6130
rect 61630 6078 61682 6130
rect 62862 6078 62914 6130
rect 65550 6078 65602 6130
rect 66558 6078 66610 6130
rect 67678 6078 67730 6130
rect 67790 6078 67842 6130
rect 69470 6078 69522 6130
rect 74734 6078 74786 6130
rect 77758 6078 77810 6130
rect 79886 6078 79938 6130
rect 81454 6078 81506 6130
rect 81678 6078 81730 6130
rect 82350 6078 82402 6130
rect 82574 6078 82626 6130
rect 89182 6078 89234 6130
rect 90750 6078 90802 6130
rect 93102 6078 93154 6130
rect 93662 6078 93714 6130
rect 95006 6078 95058 6130
rect 96126 6078 96178 6130
rect 99262 6078 99314 6130
rect 100718 6078 100770 6130
rect 101726 6078 101778 6130
rect 103070 6078 103122 6130
rect 114046 6078 114098 6130
rect 114382 6078 114434 6130
rect 116062 6078 116114 6130
rect 116958 6078 117010 6130
rect 127262 6078 127314 6130
rect 128046 6078 128098 6130
rect 133870 6078 133922 6130
rect 134654 6078 134706 6130
rect 136222 6078 136274 6130
rect 137006 6078 137058 6130
rect 139918 6078 139970 6130
rect 140814 6078 140866 6130
rect 142494 6078 142546 6130
rect 8430 5966 8482 6018
rect 13470 5966 13522 6018
rect 14366 5966 14418 6018
rect 14926 5966 14978 6018
rect 15038 5966 15090 6018
rect 18398 5966 18450 6018
rect 18958 5966 19010 6018
rect 20302 5966 20354 6018
rect 21534 5966 21586 6018
rect 26462 5966 26514 6018
rect 34190 5966 34242 6018
rect 37774 5966 37826 6018
rect 39230 5966 39282 6018
rect 40462 5966 40514 6018
rect 40798 5966 40850 6018
rect 42478 5966 42530 6018
rect 42702 5966 42754 6018
rect 44158 5966 44210 6018
rect 44606 5966 44658 6018
rect 44830 5966 44882 6018
rect 47630 5966 47682 6018
rect 48862 5966 48914 6018
rect 52222 5966 52274 6018
rect 55694 5966 55746 6018
rect 57486 5966 57538 6018
rect 57710 5966 57762 6018
rect 58046 5966 58098 6018
rect 60734 5966 60786 6018
rect 61294 5966 61346 6018
rect 61518 5966 61570 6018
rect 61854 5966 61906 6018
rect 63422 5966 63474 6018
rect 63646 5966 63698 6018
rect 64318 5966 64370 6018
rect 64654 5966 64706 6018
rect 66110 5966 66162 6018
rect 66334 5966 66386 6018
rect 67230 5966 67282 6018
rect 69358 5966 69410 6018
rect 74062 5966 74114 6018
rect 75182 5966 75234 6018
rect 77646 5966 77698 6018
rect 79102 5966 79154 6018
rect 80446 5966 80498 6018
rect 81342 5966 81394 6018
rect 84030 5966 84082 6018
rect 86046 5966 86098 6018
rect 87838 5966 87890 6018
rect 88174 5966 88226 6018
rect 90414 5966 90466 6018
rect 91646 5966 91698 6018
rect 91870 5966 91922 6018
rect 92542 5966 92594 6018
rect 92654 5966 92706 6018
rect 95566 5966 95618 6018
rect 96238 5966 96290 6018
rect 99822 5966 99874 6018
rect 100158 5966 100210 6018
rect 101838 5966 101890 6018
rect 102958 5966 103010 6018
rect 104078 5966 104130 6018
rect 104414 5966 104466 6018
rect 106878 5966 106930 6018
rect 107102 5966 107154 6018
rect 107998 5966 108050 6018
rect 108334 5966 108386 6018
rect 115278 5966 115330 6018
rect 115614 5966 115666 6018
rect 117630 5966 117682 6018
rect 121214 5966 121266 6018
rect 123118 5966 123170 6018
rect 123790 5966 123842 6018
rect 124910 5966 124962 6018
rect 129054 5966 129106 6018
rect 130846 5966 130898 6018
rect 131182 5966 131234 6018
rect 131742 5966 131794 6018
rect 132638 5966 132690 6018
rect 132974 5966 133026 6018
rect 133758 5966 133810 6018
rect 134542 5966 134594 6018
rect 135774 5966 135826 6018
rect 138350 5966 138402 6018
rect 140702 5966 140754 6018
rect 141710 5966 141762 6018
rect 142382 5966 142434 6018
rect 143390 5966 143442 6018
rect 145294 5966 145346 6018
rect 146750 5966 146802 6018
rect 8654 5854 8706 5906
rect 13246 5854 13298 5906
rect 14030 5854 14082 5906
rect 15710 5854 15762 5906
rect 16606 5854 16658 5906
rect 20638 5854 20690 5906
rect 21198 5854 21250 5906
rect 22430 5854 22482 5906
rect 24110 5854 24162 5906
rect 25678 5854 25730 5906
rect 30942 5854 30994 5906
rect 32622 5854 32674 5906
rect 33854 5854 33906 5906
rect 34750 5854 34802 5906
rect 38558 5854 38610 5906
rect 39454 5854 39506 5906
rect 42366 5854 42418 5906
rect 42926 5854 42978 5906
rect 45278 5854 45330 5906
rect 46622 5854 46674 5906
rect 47406 5854 47458 5906
rect 47966 5854 48018 5906
rect 49982 5854 50034 5906
rect 55470 5854 55522 5906
rect 56254 5854 56306 5906
rect 58942 5854 58994 5906
rect 59614 5854 59666 5906
rect 60398 5854 60450 5906
rect 62526 5854 62578 5906
rect 66782 5854 66834 5906
rect 67454 5854 67506 5906
rect 67566 5854 67618 5906
rect 68462 5854 68514 5906
rect 68798 5854 68850 5906
rect 69134 5854 69186 5906
rect 70030 5854 70082 5906
rect 70254 5854 70306 5906
rect 71934 5854 71986 5906
rect 72606 5854 72658 5906
rect 73390 5854 73442 5906
rect 73614 5854 73666 5906
rect 73950 5854 74002 5906
rect 74398 5854 74450 5906
rect 75406 5854 75458 5906
rect 76526 5854 76578 5906
rect 77982 5854 78034 5906
rect 78094 5854 78146 5906
rect 78878 5854 78930 5906
rect 80334 5854 80386 5906
rect 80670 5854 80722 5906
rect 82126 5854 82178 5906
rect 82686 5854 82738 5906
rect 83470 5854 83522 5906
rect 85486 5854 85538 5906
rect 89742 5854 89794 5906
rect 89966 5854 90018 5906
rect 90078 5854 90130 5906
rect 90750 5854 90802 5906
rect 94670 5854 94722 5906
rect 96462 5854 96514 5906
rect 97470 5854 97522 5906
rect 98142 5854 98194 5906
rect 98926 5854 98978 5906
rect 101278 5854 101330 5906
rect 102062 5854 102114 5906
rect 105646 5854 105698 5906
rect 107438 5854 107490 5906
rect 109230 5854 109282 5906
rect 113150 5854 113202 5906
rect 113374 5854 113426 5906
rect 118414 5854 118466 5906
rect 119758 5854 119810 5906
rect 119870 5854 119922 5906
rect 122334 5854 122386 5906
rect 124126 5854 124178 5906
rect 128270 5854 128322 5906
rect 129278 5854 129330 5906
rect 130286 5854 130338 5906
rect 134878 5854 134930 5906
rect 135438 5854 135490 5906
rect 137342 5854 137394 5906
rect 140142 5854 140194 5906
rect 141038 5854 141090 5906
rect 142718 5854 142770 5906
rect 145518 5854 145570 5906
rect 7982 5742 8034 5794
rect 9662 5742 9714 5794
rect 11230 5742 11282 5794
rect 11790 5742 11842 5794
rect 12686 5742 12738 5794
rect 19854 5742 19906 5794
rect 28590 5742 28642 5794
rect 29934 5742 29986 5794
rect 31614 5742 31666 5794
rect 32062 5742 32114 5794
rect 35086 5742 35138 5794
rect 35646 5742 35698 5794
rect 40014 5742 40066 5794
rect 45054 5742 45106 5794
rect 57934 5742 57986 5794
rect 58606 5742 58658 5794
rect 59502 5742 59554 5794
rect 63758 5742 63810 5794
rect 65438 5742 65490 5794
rect 70926 5742 70978 5794
rect 71822 5742 71874 5794
rect 74734 5742 74786 5794
rect 76190 5742 76242 5794
rect 77086 5742 77138 5794
rect 82462 5742 82514 5794
rect 85598 5742 85650 5794
rect 90974 5742 91026 5794
rect 91758 5742 91810 5794
rect 93998 5742 94050 5794
rect 95790 5742 95842 5794
rect 105422 5742 105474 5794
rect 106318 5742 106370 5794
rect 107326 5742 107378 5794
rect 109902 5742 109954 5794
rect 112142 5742 112194 5794
rect 113598 5742 113650 5794
rect 116510 5742 116562 5794
rect 121102 5742 121154 5794
rect 121438 5742 121490 5794
rect 121998 5742 122050 5794
rect 122110 5742 122162 5794
rect 124014 5742 124066 5794
rect 125582 5742 125634 5794
rect 126030 5742 126082 5794
rect 126478 5742 126530 5794
rect 126814 5742 126866 5794
rect 137790 5742 137842 5794
rect 138910 5742 138962 5794
rect 143950 5742 144002 5794
rect 146078 5742 146130 5794
rect 147310 5742 147362 5794
rect 147758 5742 147810 5794
rect 148206 5742 148258 5794
rect 148766 5742 148818 5794
rect 149102 5742 149154 5794
rect 149662 5742 149714 5794
rect 149998 5742 150050 5794
rect 17838 5630 17890 5682
rect 18174 5630 18226 5682
rect 28926 5630 28978 5682
rect 29486 5630 29538 5682
rect 43374 5630 43426 5682
rect 68910 5630 68962 5682
rect 92542 5630 92594 5682
rect 93326 5630 93378 5682
rect 93998 5630 94050 5682
rect 96014 5630 96066 5682
rect 97358 5630 97410 5682
rect 101502 5630 101554 5682
rect 103070 5630 103122 5682
rect 117742 5630 117794 5682
rect 118526 5630 118578 5682
rect 118750 5630 118802 5682
rect 118862 5630 118914 5682
rect 119422 5630 119474 5682
rect 119534 5630 119586 5682
rect 126030 5630 126082 5682
rect 126254 5630 126306 5682
rect 126478 5630 126530 5682
rect 126702 5630 126754 5682
rect 127038 5630 127090 5682
rect 127374 5630 127426 5682
rect 127934 5630 127986 5682
rect 129950 5630 130002 5682
rect 130286 5630 130338 5682
rect 133982 5630 134034 5682
rect 139806 5630 139858 5682
rect 148654 5630 148706 5682
rect 149102 5630 149154 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 96638 5462 96690 5514
rect 96742 5462 96794 5514
rect 96846 5462 96898 5514
rect 127358 5462 127410 5514
rect 127462 5462 127514 5514
rect 127566 5462 127618 5514
rect 158078 5462 158130 5514
rect 158182 5462 158234 5514
rect 158286 5462 158338 5514
rect 8990 5294 9042 5346
rect 14590 5294 14642 5346
rect 45950 5294 46002 5346
rect 46286 5294 46338 5346
rect 62302 5294 62354 5346
rect 62638 5294 62690 5346
rect 68462 5294 68514 5346
rect 69806 5294 69858 5346
rect 71374 5294 71426 5346
rect 79998 5294 80050 5346
rect 80894 5294 80946 5346
rect 95902 5294 95954 5346
rect 96238 5294 96290 5346
rect 102062 5294 102114 5346
rect 106766 5294 106818 5346
rect 106990 5294 107042 5346
rect 110238 5294 110290 5346
rect 111134 5294 111186 5346
rect 111470 5294 111522 5346
rect 119646 5294 119698 5346
rect 123006 5294 123058 5346
rect 123454 5294 123506 5346
rect 123902 5294 123954 5346
rect 125582 5294 125634 5346
rect 125806 5294 125858 5346
rect 133086 5294 133138 5346
rect 133198 5294 133250 5346
rect 133422 5294 133474 5346
rect 136670 5294 136722 5346
rect 136782 5294 136834 5346
rect 137006 5294 137058 5346
rect 137230 5294 137282 5346
rect 139134 5294 139186 5346
rect 139694 5294 139746 5346
rect 8430 5182 8482 5234
rect 13694 5182 13746 5234
rect 18958 5182 19010 5234
rect 19854 5182 19906 5234
rect 21870 5182 21922 5234
rect 24110 5182 24162 5234
rect 27806 5182 27858 5234
rect 30718 5182 30770 5234
rect 31502 5182 31554 5234
rect 33070 5182 33122 5234
rect 36878 5182 36930 5234
rect 40462 5182 40514 5234
rect 42590 5182 42642 5234
rect 47406 5182 47458 5234
rect 49758 5182 49810 5234
rect 51886 5182 51938 5234
rect 54574 5182 54626 5234
rect 56702 5182 56754 5234
rect 58494 5182 58546 5234
rect 60622 5182 60674 5234
rect 68238 5182 68290 5234
rect 70030 5182 70082 5234
rect 75294 5182 75346 5234
rect 75630 5182 75682 5234
rect 78206 5182 78258 5234
rect 78654 5182 78706 5234
rect 81230 5182 81282 5234
rect 84254 5182 84306 5234
rect 87390 5182 87442 5234
rect 87502 5182 87554 5234
rect 87614 5182 87666 5234
rect 88174 5182 88226 5234
rect 88958 5182 89010 5234
rect 91310 5182 91362 5234
rect 91646 5182 91698 5234
rect 97806 5182 97858 5234
rect 98030 5182 98082 5234
rect 99598 5182 99650 5234
rect 99822 5182 99874 5234
rect 100270 5182 100322 5234
rect 101054 5182 101106 5234
rect 102286 5182 102338 5234
rect 106318 5182 106370 5234
rect 106654 5182 106706 5234
rect 107774 5182 107826 5234
rect 112254 5182 112306 5234
rect 113822 5182 113874 5234
rect 119870 5182 119922 5234
rect 119982 5182 120034 5234
rect 121662 5182 121714 5234
rect 121774 5182 121826 5234
rect 121886 5182 121938 5234
rect 126030 5182 126082 5234
rect 131742 5182 131794 5234
rect 137790 5182 137842 5234
rect 7646 5070 7698 5122
rect 8654 5070 8706 5122
rect 12014 5070 12066 5122
rect 14254 5070 14306 5122
rect 16158 5070 16210 5122
rect 16830 5070 16882 5122
rect 20750 5070 20802 5122
rect 23438 5070 23490 5122
rect 26910 5070 26962 5122
rect 28702 5070 28754 5122
rect 32286 5070 32338 5122
rect 35982 5070 36034 5122
rect 37886 5070 37938 5122
rect 38222 5070 38274 5122
rect 43262 5070 43314 5122
rect 43934 5070 43986 5122
rect 45390 5070 45442 5122
rect 48078 5070 48130 5122
rect 52558 5070 52610 5122
rect 53790 5070 53842 5122
rect 57710 5070 57762 5122
rect 61854 5070 61906 5122
rect 66334 5070 66386 5122
rect 66782 5070 66834 5122
rect 67678 5070 67730 5122
rect 70254 5070 70306 5122
rect 72270 5070 72322 5122
rect 73614 5070 73666 5122
rect 77646 5070 77698 5122
rect 81902 5070 81954 5122
rect 83582 5070 83634 5122
rect 84478 5070 84530 5122
rect 85486 5070 85538 5122
rect 86718 5070 86770 5122
rect 87166 5070 87218 5122
rect 89070 5070 89122 5122
rect 90638 5070 90690 5122
rect 97134 5070 97186 5122
rect 98590 5070 98642 5122
rect 98926 5070 98978 5122
rect 101614 5070 101666 5122
rect 102510 5070 102562 5122
rect 103742 5070 103794 5122
rect 104190 5070 104242 5122
rect 105310 5070 105362 5122
rect 105646 5070 105698 5122
rect 107662 5070 107714 5122
rect 109454 5070 109506 5122
rect 110238 5070 110290 5122
rect 112590 5070 112642 5122
rect 113934 5070 113986 5122
rect 115278 5070 115330 5122
rect 119198 5070 119250 5122
rect 120094 5070 120146 5122
rect 121214 5070 121266 5122
rect 123678 5070 123730 5122
rect 124910 5070 124962 5122
rect 125358 5070 125410 5122
rect 127262 5070 127314 5122
rect 127710 5070 127762 5122
rect 127934 5070 127986 5122
rect 128158 5070 128210 5122
rect 128382 5070 128434 5122
rect 128942 5070 128994 5122
rect 130510 5070 130562 5122
rect 130734 5070 130786 5122
rect 133646 5070 133698 5122
rect 142942 5294 142994 5346
rect 143950 5294 144002 5346
rect 147646 5182 147698 5234
rect 135998 5070 136050 5122
rect 139806 5070 139858 5122
rect 143054 5070 143106 5122
rect 143278 5070 143330 5122
rect 144062 5070 144114 5122
rect 149102 5070 149154 5122
rect 152462 5070 152514 5122
rect 159294 5070 159346 5122
rect 161086 5070 161138 5122
rect 7870 4958 7922 5010
rect 9550 4958 9602 5010
rect 9886 4958 9938 5010
rect 11230 4958 11282 5010
rect 11566 4958 11618 5010
rect 12910 4958 12962 5010
rect 14814 4958 14866 5010
rect 15150 4958 15202 5010
rect 22654 4958 22706 5010
rect 26238 4958 26290 5010
rect 30270 4958 30322 5010
rect 35198 4958 35250 5010
rect 37550 4958 37602 5010
rect 37998 4958 38050 5010
rect 38670 4958 38722 5010
rect 39006 4958 39058 5010
rect 39566 4958 39618 5010
rect 44382 4958 44434 5010
rect 44718 4958 44770 5010
rect 48862 4958 48914 5010
rect 49198 4958 49250 5010
rect 61518 4958 61570 5010
rect 64094 4958 64146 5010
rect 64430 4958 64482 5010
rect 64990 4958 65042 5010
rect 65326 4958 65378 5010
rect 66894 4958 66946 5010
rect 69358 4958 69410 5010
rect 69582 4958 69634 5010
rect 70814 4958 70866 5010
rect 71038 4958 71090 5010
rect 71262 4958 71314 5010
rect 72494 4958 72546 5010
rect 73502 4958 73554 5010
rect 76190 4958 76242 5010
rect 77982 4958 78034 5010
rect 79102 4958 79154 5010
rect 79438 4958 79490 5010
rect 80222 4958 80274 5010
rect 81118 4958 81170 5010
rect 83470 4958 83522 5010
rect 83918 4958 83970 5010
rect 86494 4958 86546 5010
rect 89742 4958 89794 5010
rect 90414 4958 90466 5010
rect 90974 4958 91026 5010
rect 91422 4958 91474 5010
rect 92430 4958 92482 5010
rect 93214 4958 93266 5010
rect 94110 4958 94162 5010
rect 95006 4958 95058 5010
rect 96126 4958 96178 5010
rect 96910 4958 96962 5010
rect 97470 4958 97522 5010
rect 98814 4958 98866 5010
rect 99262 4958 99314 5010
rect 101838 4958 101890 5010
rect 102398 4958 102450 5010
rect 103070 4958 103122 5010
rect 104750 4958 104802 5010
rect 105982 4958 106034 5010
rect 108334 4958 108386 5010
rect 110574 4958 110626 5010
rect 113038 4958 113090 5010
rect 114606 4958 114658 5010
rect 117070 4958 117122 5010
rect 117406 4958 117458 5010
rect 118302 4958 118354 5010
rect 118638 4958 118690 5010
rect 119422 4958 119474 5010
rect 120766 4958 120818 5010
rect 121326 4958 121378 5010
rect 124126 4958 124178 5010
rect 129278 4958 129330 5010
rect 130622 4958 130674 5010
rect 131070 4958 131122 5010
rect 131630 4958 131682 5010
rect 133758 4958 133810 5010
rect 134318 4958 134370 5010
rect 134654 4958 134706 5010
rect 135438 4958 135490 5010
rect 135662 4958 135714 5010
rect 137342 4958 137394 5010
rect 137902 4958 137954 5010
rect 138350 4958 138402 5010
rect 138574 4958 138626 5010
rect 139358 4958 139410 5010
rect 140926 4958 140978 5010
rect 141262 4958 141314 5010
rect 141822 4958 141874 5010
rect 142158 4958 142210 5010
rect 143390 4958 143442 5010
rect 144958 4958 145010 5010
rect 145294 4958 145346 5010
rect 146190 4958 146242 5010
rect 146750 4958 146802 5010
rect 147086 4958 147138 5010
rect 147758 4958 147810 5010
rect 148878 4958 148930 5010
rect 7086 4846 7138 4898
rect 10782 4846 10834 4898
rect 12574 4846 12626 4898
rect 29934 4846 29986 4898
rect 39902 4846 39954 4898
rect 46174 4846 46226 4898
rect 57262 4846 57314 4898
rect 63646 4846 63698 4898
rect 69694 4846 69746 4898
rect 76526 4846 76578 4898
rect 77422 4846 77474 4898
rect 77534 4846 77586 4898
rect 78094 4846 78146 4898
rect 80110 4846 80162 4898
rect 82126 4846 82178 4898
rect 82686 4846 82738 4898
rect 83358 4846 83410 4898
rect 84030 4846 84082 4898
rect 85822 4846 85874 4898
rect 86606 4846 86658 4898
rect 90526 4846 90578 4898
rect 92094 4846 92146 4898
rect 93550 4846 93602 4898
rect 94446 4846 94498 4898
rect 95342 4846 95394 4898
rect 97022 4846 97074 4898
rect 97582 4846 97634 4898
rect 99374 4846 99426 4898
rect 103630 4846 103682 4898
rect 105534 4846 105586 4898
rect 106094 4846 106146 4898
rect 109118 4846 109170 4898
rect 111358 4846 111410 4898
rect 115502 4846 115554 4898
rect 115950 4846 116002 4898
rect 120878 4846 120930 4898
rect 122446 4846 122498 4898
rect 126590 4846 126642 4898
rect 129838 4846 129890 4898
rect 131854 4846 131906 4898
rect 135886 4846 135938 4898
rect 138126 4846 138178 4898
rect 139246 4846 139298 4898
rect 140030 4846 140082 4898
rect 144174 4846 144226 4898
rect 145854 4846 145906 4898
rect 147870 4846 147922 4898
rect 150110 4846 150162 4898
rect 150670 4846 150722 4898
rect 151230 4846 151282 4898
rect 151790 4846 151842 4898
rect 155374 4846 155426 4898
rect 156718 4846 156770 4898
rect 158398 4846 158450 4898
rect 161534 4846 161586 4898
rect 167134 4846 167186 4898
rect 168030 4846 168082 4898
rect 168926 4846 168978 4898
rect 169374 4846 169426 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 81278 4678 81330 4730
rect 81382 4678 81434 4730
rect 81486 4678 81538 4730
rect 111998 4678 112050 4730
rect 112102 4678 112154 4730
rect 112206 4678 112258 4730
rect 142718 4678 142770 4730
rect 142822 4678 142874 4730
rect 142926 4678 142978 4730
rect 173438 4678 173490 4730
rect 173542 4678 173594 4730
rect 173646 4678 173698 4730
rect 10446 4510 10498 4562
rect 16046 4510 16098 4562
rect 16606 4510 16658 4562
rect 18734 4510 18786 4562
rect 23102 4510 23154 4562
rect 26014 4510 26066 4562
rect 26686 4510 26738 4562
rect 33518 4510 33570 4562
rect 39454 4510 39506 4562
rect 40574 4510 40626 4562
rect 40798 4510 40850 4562
rect 57822 4510 57874 4562
rect 61854 4510 61906 4562
rect 62638 4510 62690 4562
rect 64318 4510 64370 4562
rect 67790 4510 67842 4562
rect 68910 4510 68962 4562
rect 71374 4510 71426 4562
rect 72158 4510 72210 4562
rect 74174 4510 74226 4562
rect 78542 4510 78594 4562
rect 78654 4510 78706 4562
rect 81566 4510 81618 4562
rect 83694 4510 83746 4562
rect 84478 4510 84530 4562
rect 84590 4510 84642 4562
rect 85150 4510 85202 4562
rect 90078 4510 90130 4562
rect 90190 4510 90242 4562
rect 91086 4510 91138 4562
rect 93326 4510 93378 4562
rect 96350 4510 96402 4562
rect 100158 4510 100210 4562
rect 100270 4510 100322 4562
rect 100382 4510 100434 4562
rect 101054 4510 101106 4562
rect 102062 4510 102114 4562
rect 105310 4510 105362 4562
rect 105422 4510 105474 4562
rect 108334 4510 108386 4562
rect 109230 4510 109282 4562
rect 113262 4510 113314 4562
rect 113374 4510 113426 4562
rect 113934 4510 113986 4562
rect 114942 4510 114994 4562
rect 115726 4510 115778 4562
rect 116846 4510 116898 4562
rect 117406 4510 117458 4562
rect 117518 4510 117570 4562
rect 118078 4510 118130 4562
rect 119758 4510 119810 4562
rect 121326 4510 121378 4562
rect 122222 4510 122274 4562
rect 122782 4510 122834 4562
rect 123454 4510 123506 4562
rect 123678 4510 123730 4562
rect 124574 4510 124626 4562
rect 126366 4510 126418 4562
rect 127934 4510 127986 4562
rect 133758 4510 133810 4562
rect 135326 4510 135378 4562
rect 138238 4510 138290 4562
rect 139694 4510 139746 4562
rect 141374 4510 141426 4562
rect 141710 4510 141762 4562
rect 11454 4398 11506 4450
rect 12798 4398 12850 4450
rect 20078 4398 20130 4450
rect 27582 4398 27634 4450
rect 29934 4398 29986 4450
rect 37998 4398 38050 4450
rect 39342 4398 39394 4450
rect 40126 4398 40178 4450
rect 42366 4398 42418 4450
rect 43262 4398 43314 4450
rect 47630 4398 47682 4450
rect 51998 4398 52050 4450
rect 60510 4398 60562 4450
rect 62302 4398 62354 4450
rect 63198 4398 63250 4450
rect 63534 4398 63586 4450
rect 64430 4398 64482 4450
rect 67678 4398 67730 4450
rect 68350 4398 68402 4450
rect 71822 4398 71874 4450
rect 74062 4398 74114 4450
rect 75630 4398 75682 4450
rect 78430 4398 78482 4450
rect 82014 4398 82066 4450
rect 82350 4398 82402 4450
rect 85038 4398 85090 4450
rect 86382 4398 86434 4450
rect 86718 4398 86770 4450
rect 89294 4398 89346 4450
rect 90638 4398 90690 4450
rect 92094 4398 92146 4450
rect 97358 4398 97410 4450
rect 97470 4398 97522 4450
rect 99822 4398 99874 4450
rect 102958 4398 103010 4450
rect 103294 4398 103346 4450
rect 104414 4398 104466 4450
rect 108894 4398 108946 4450
rect 112030 4398 112082 4450
rect 112366 4398 112418 4450
rect 113822 4398 113874 4450
rect 116174 4398 116226 4450
rect 117966 4398 118018 4450
rect 119422 4398 119474 4450
rect 119646 4398 119698 4450
rect 120318 4398 120370 4450
rect 121774 4398 121826 4450
rect 125582 4398 125634 4450
rect 125806 4398 125858 4450
rect 127822 4398 127874 4450
rect 129054 4398 129106 4450
rect 129278 4398 129330 4450
rect 130062 4398 130114 4450
rect 130286 4398 130338 4450
rect 130846 4398 130898 4450
rect 131070 4398 131122 4450
rect 131742 4398 131794 4450
rect 131966 4398 132018 4450
rect 132974 4398 133026 4450
rect 133198 4398 133250 4450
rect 133422 4398 133474 4450
rect 133870 4398 133922 4450
rect 134766 4398 134818 4450
rect 135662 4398 135714 4450
rect 136110 4398 136162 4450
rect 137006 4398 137058 4450
rect 139582 4398 139634 4450
rect 139806 4398 139858 4450
rect 140366 4398 140418 4450
rect 8542 4286 8594 4338
rect 10110 4286 10162 4338
rect 11230 4286 11282 4338
rect 12126 4286 12178 4338
rect 15822 4286 15874 4338
rect 16942 4286 16994 4338
rect 18398 4286 18450 4338
rect 19294 4286 19346 4338
rect 22878 4286 22930 4338
rect 23774 4286 23826 4338
rect 25790 4286 25842 4338
rect 27022 4286 27074 4338
rect 27470 4286 27522 4338
rect 29150 4286 29202 4338
rect 32846 4286 32898 4338
rect 34302 4286 34354 4338
rect 38670 4286 38722 4338
rect 39678 4286 39730 4338
rect 40350 4286 40402 4338
rect 40798 4286 40850 4338
rect 42254 4286 42306 4338
rect 42590 4286 42642 4338
rect 42814 4286 42866 4338
rect 44942 4286 44994 4338
rect 48414 4286 48466 4338
rect 53902 4286 53954 4338
rect 56590 4286 56642 4338
rect 57486 4286 57538 4338
rect 61182 4286 61234 4338
rect 64094 4286 64146 4338
rect 65550 4286 65602 4338
rect 67342 4286 67394 4338
rect 67902 4286 67954 4338
rect 68126 4286 68178 4338
rect 69358 4286 69410 4338
rect 71150 4286 71202 4338
rect 71710 4286 71762 4338
rect 72382 4286 72434 4338
rect 73390 4286 73442 4338
rect 73614 4286 73666 4338
rect 73726 4286 73778 4338
rect 74398 4286 74450 4338
rect 75406 4286 75458 4338
rect 76190 4286 76242 4338
rect 79326 4286 79378 4338
rect 82798 4286 82850 4338
rect 83246 4286 83298 4338
rect 83358 4286 83410 4338
rect 83582 4286 83634 4338
rect 83806 4286 83858 4338
rect 84702 4286 84754 4338
rect 85374 4286 85426 4338
rect 85598 4286 85650 4338
rect 88286 4286 88338 4338
rect 89406 4286 89458 4338
rect 90302 4286 90354 4338
rect 91198 4286 91250 4338
rect 91758 4286 91810 4338
rect 92766 4286 92818 4338
rect 92990 4286 93042 4338
rect 94670 4286 94722 4338
rect 98254 4286 98306 4338
rect 100046 4286 100098 4338
rect 101166 4286 101218 4338
rect 101726 4286 101778 4338
rect 101950 4286 102002 4338
rect 102174 4286 102226 4338
rect 102398 4286 102450 4338
rect 104190 4286 104242 4338
rect 105646 4286 105698 4338
rect 105982 4286 106034 4338
rect 106542 4286 106594 4338
rect 108446 4286 108498 4338
rect 108558 4286 108610 4338
rect 109230 4286 109282 4338
rect 111022 4286 111074 4338
rect 113710 4286 113762 4338
rect 114158 4286 114210 4338
rect 115502 4286 115554 4338
rect 116062 4286 116114 4338
rect 116510 4286 116562 4338
rect 116734 4286 116786 4338
rect 117630 4286 117682 4338
rect 119870 4286 119922 4338
rect 121214 4286 121266 4338
rect 121438 4286 121490 4338
rect 122110 4286 122162 4338
rect 122334 4286 122386 4338
rect 124014 4286 124066 4338
rect 124798 4286 124850 4338
rect 126702 4286 126754 4338
rect 132638 4286 132690 4338
rect 133534 4286 133586 4338
rect 134430 4286 134482 4338
rect 137342 4286 137394 4338
rect 137566 4286 137618 4338
rect 138126 4286 138178 4338
rect 138350 4286 138402 4338
rect 138798 4286 138850 4338
rect 140590 4286 140642 4338
rect 6862 4174 6914 4226
rect 7534 4174 7586 4226
rect 9102 4174 9154 4226
rect 14926 4174 14978 4226
rect 17838 4174 17890 4226
rect 22206 4174 22258 4226
rect 24446 4174 24498 4226
rect 28590 4174 28642 4226
rect 32062 4174 32114 4226
rect 34750 4174 34802 4226
rect 35870 4174 35922 4226
rect 41694 4174 41746 4226
rect 44270 4174 44322 4226
rect 45502 4174 45554 4226
rect 55582 4174 55634 4226
rect 58382 4174 58434 4226
rect 66110 4174 66162 4226
rect 70030 4174 70082 4226
rect 72046 4174 72098 4226
rect 74622 4174 74674 4226
rect 76862 4174 76914 4226
rect 77982 4174 78034 4226
rect 79998 4174 80050 4226
rect 87726 4174 87778 4226
rect 90974 4174 91026 4226
rect 93774 4174 93826 4226
rect 95342 4174 95394 4226
rect 98702 4174 98754 4226
rect 107102 4174 107154 4226
rect 109454 4174 109506 4226
rect 110238 4174 110290 4226
rect 114494 4174 114546 4226
rect 118190 4174 118242 4226
rect 118638 4174 118690 4226
rect 120094 4174 120146 4226
rect 123566 4174 123618 4226
rect 125470 4174 125522 4226
rect 127150 4174 127202 4226
rect 129166 4174 129218 4226
rect 129950 4174 130002 4226
rect 131182 4174 131234 4226
rect 132078 4174 132130 4226
rect 134542 4174 134594 4226
rect 137118 4174 137170 4226
rect 128046 4062 128098 4114
rect 144062 4510 144114 4562
rect 146078 4510 146130 4562
rect 151230 4510 151282 4562
rect 156270 4510 156322 4562
rect 159070 4510 159122 4562
rect 161310 4510 161362 4562
rect 144958 4398 145010 4450
rect 145518 4398 145570 4450
rect 146974 4398 147026 4450
rect 147870 4398 147922 4450
rect 148094 4398 148146 4450
rect 149662 4398 149714 4450
rect 149998 4398 150050 4450
rect 150558 4398 150610 4450
rect 153470 4398 153522 4450
rect 155150 4398 155202 4450
rect 157166 4398 157218 4450
rect 158398 4398 158450 4450
rect 159966 4398 160018 4450
rect 162206 4398 162258 4450
rect 163550 4398 163602 4450
rect 165230 4398 165282 4450
rect 166910 4398 166962 4450
rect 168030 4398 168082 4450
rect 169150 4398 169202 4450
rect 170270 4398 170322 4450
rect 171950 4398 172002 4450
rect 173070 4398 173122 4450
rect 141598 4286 141650 4338
rect 141822 4286 141874 4338
rect 142046 4286 142098 4338
rect 142830 4286 142882 4338
rect 143278 4286 143330 4338
rect 143502 4286 143554 4338
rect 145070 4286 145122 4338
rect 145182 4286 145234 4338
rect 146302 4286 146354 4338
rect 147310 4286 147362 4338
rect 148766 4286 148818 4338
rect 149102 4286 149154 4338
rect 151454 4286 151506 4338
rect 156494 4286 156546 4338
rect 161534 4286 161586 4338
rect 169374 4286 169426 4338
rect 142270 4174 142322 4226
rect 143054 4174 143106 4226
rect 144174 4174 144226 4226
rect 148990 4174 149042 4226
rect 152014 4174 152066 4226
rect 152798 4174 152850 4226
rect 154030 4174 154082 4226
rect 154590 4174 154642 4226
rect 155822 4174 155874 4226
rect 157726 4174 157778 4226
rect 159182 4174 159234 4226
rect 160750 4174 160802 4226
rect 162766 4174 162818 4226
rect 164110 4174 164162 4226
rect 164558 4174 164610 4226
rect 165790 4174 165842 4226
rect 166350 4174 166402 4226
rect 170830 4174 170882 4226
rect 171390 4174 171442 4226
rect 172510 4174 172562 4226
rect 173630 4174 173682 4226
rect 138574 4062 138626 4114
rect 141374 4062 141426 4114
rect 147310 4062 147362 4114
rect 148206 4062 148258 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 96638 3894 96690 3946
rect 96742 3894 96794 3946
rect 96846 3894 96898 3946
rect 127358 3894 127410 3946
rect 127462 3894 127514 3946
rect 127566 3894 127618 3946
rect 158078 3894 158130 3946
rect 158182 3894 158234 3946
rect 158286 3894 158338 3946
rect 21534 3726 21586 3778
rect 21870 3726 21922 3778
rect 26350 3726 26402 3778
rect 26686 3726 26738 3778
rect 30382 3726 30434 3778
rect 30718 3726 30770 3778
rect 64318 3726 64370 3778
rect 64990 3726 65042 3778
rect 76974 3726 77026 3778
rect 8318 3614 8370 3666
rect 10334 3614 10386 3666
rect 12574 3614 12626 3666
rect 13806 3614 13858 3666
rect 32510 3614 32562 3666
rect 37886 3614 37938 3666
rect 39566 3614 39618 3666
rect 41806 3614 41858 3666
rect 43150 3614 43202 3666
rect 49086 3614 49138 3666
rect 51214 3614 51266 3666
rect 53118 3614 53170 3666
rect 61406 3614 61458 3666
rect 63086 3614 63138 3666
rect 64766 3614 64818 3666
rect 71038 3614 71090 3666
rect 72718 3614 72770 3666
rect 76526 3614 76578 3666
rect 77086 3614 77138 3666
rect 81006 3614 81058 3666
rect 82798 3614 82850 3666
rect 86270 3614 86322 3666
rect 88286 3614 88338 3666
rect 88734 3614 88786 3666
rect 89182 3614 89234 3666
rect 95790 3614 95842 3666
rect 98926 3614 98978 3666
rect 104974 3614 105026 3666
rect 105534 3614 105586 3666
rect 109902 3614 109954 3666
rect 110350 3614 110402 3666
rect 114046 3614 114098 3666
rect 117966 3614 118018 3666
rect 121774 3614 121826 3666
rect 129950 3614 130002 3666
rect 148766 3614 148818 3666
rect 6526 3502 6578 3554
rect 10782 3502 10834 3554
rect 11678 3502 11730 3554
rect 14254 3502 14306 3554
rect 15150 3502 15202 3554
rect 18734 3502 18786 3554
rect 20638 3502 20690 3554
rect 22542 3502 22594 3554
rect 24558 3502 24610 3554
rect 25454 3502 25506 3554
rect 27470 3502 27522 3554
rect 28254 3502 28306 3554
rect 29486 3502 29538 3554
rect 34414 3502 34466 3554
rect 36318 3502 36370 3554
rect 37438 3502 37490 3554
rect 40238 3502 40290 3554
rect 41134 3502 41186 3554
rect 44046 3502 44098 3554
rect 46062 3502 46114 3554
rect 46846 3502 46898 3554
rect 51998 3502 52050 3554
rect 54126 3502 54178 3554
rect 55694 3502 55746 3554
rect 57934 3502 57986 3554
rect 59838 3502 59890 3554
rect 60846 3502 60898 3554
rect 63534 3502 63586 3554
rect 65214 3502 65266 3554
rect 66110 3502 66162 3554
rect 68462 3502 68514 3554
rect 70366 3502 70418 3554
rect 73726 3502 73778 3554
rect 74286 3502 74338 3554
rect 77310 3502 77362 3554
rect 77870 3502 77922 3554
rect 80334 3502 80386 3554
rect 82126 3502 82178 3554
rect 84254 3502 84306 3554
rect 87054 3502 87106 3554
rect 89630 3502 89682 3554
rect 92094 3502 92146 3554
rect 93774 3502 93826 3554
rect 94670 3502 94722 3554
rect 96462 3502 96514 3554
rect 98478 3502 98530 3554
rect 99934 3502 99986 3554
rect 102846 3502 102898 3554
rect 104750 3502 104802 3554
rect 105534 3502 105586 3554
rect 107550 3502 107602 3554
rect 108222 3502 108274 3554
rect 110798 3502 110850 3554
rect 112814 3502 112866 3554
rect 113374 3502 113426 3554
rect 115726 3502 115778 3554
rect 117294 3502 117346 3554
rect 119422 3502 119474 3554
rect 121214 3502 121266 3554
rect 121438 3502 121490 3554
rect 121662 3502 121714 3554
rect 123678 3502 123730 3554
rect 124462 3502 124514 3554
rect 125358 3502 125410 3554
rect 126366 3502 126418 3554
rect 127262 3502 127314 3554
rect 128494 3502 128546 3554
rect 129054 3502 129106 3554
rect 131518 3502 131570 3554
rect 132078 3502 132130 3554
rect 134206 3502 134258 3554
rect 135438 3502 135490 3554
rect 137118 3502 137170 3554
rect 138014 3502 138066 3554
rect 139022 3502 139074 3554
rect 140254 3502 140306 3554
rect 141150 3502 141202 3554
rect 143278 3502 143330 3554
rect 144174 3502 144226 3554
rect 144958 3502 145010 3554
rect 147198 3502 147250 3554
rect 148094 3502 148146 3554
rect 148990 3502 149042 3554
rect 149886 3502 149938 3554
rect 151118 3502 151170 3554
rect 151902 3502 151954 3554
rect 153694 3502 153746 3554
rect 155822 3502 155874 3554
rect 156718 3502 156770 3554
rect 157614 3502 157666 3554
rect 158958 3502 159010 3554
rect 160638 3502 160690 3554
rect 161646 3502 161698 3554
rect 163662 3502 163714 3554
rect 165454 3502 165506 3554
rect 167582 3502 167634 3554
rect 169486 3502 169538 3554
rect 170718 3502 170770 3554
rect 172398 3502 172450 3554
rect 173406 3502 173458 3554
rect 5854 3390 5906 3442
rect 16046 3390 16098 3442
rect 17838 3390 17890 3442
rect 19742 3390 19794 3442
rect 22430 3390 22482 3442
rect 23662 3390 23714 3442
rect 27246 3390 27298 3442
rect 30942 3390 30994 3442
rect 31502 3390 31554 3442
rect 33518 3390 33570 3442
rect 35422 3390 35474 3442
rect 45390 3390 45442 3442
rect 47742 3390 47794 3442
rect 55022 3390 55074 3442
rect 57150 3390 57202 3442
rect 58942 3390 58994 3442
rect 67006 3390 67058 3442
rect 69358 3390 69410 3442
rect 75182 3390 75234 3442
rect 78766 3390 78818 3442
rect 85150 3390 85202 3442
rect 90526 3390 90578 3442
rect 92878 3390 92930 3442
rect 97246 3390 97298 3442
rect 100718 3390 100770 3442
rect 101950 3390 102002 3442
rect 104078 3390 104130 3442
rect 106430 3390 106482 3442
rect 109006 3390 109058 3442
rect 111918 3390 111970 3442
rect 116398 3390 116450 3442
rect 120318 3390 120370 3442
rect 121774 3390 121826 3442
rect 130174 3390 130226 3442
rect 133310 3390 133362 3442
rect 135102 3390 135154 3442
rect 136334 3390 136386 3442
rect 142046 3390 142098 3442
rect 145630 3390 145682 3442
rect 145966 3390 146018 3442
rect 148654 3390 148706 3442
rect 152910 3390 152962 3442
rect 155038 3390 155090 3442
rect 157390 3390 157442 3442
rect 159854 3390 159906 3442
rect 162878 3390 162930 3442
rect 164670 3390 164722 3442
rect 166798 3390 166850 3442
rect 168590 3390 168642 3442
rect 171614 3390 171666 3442
rect 14590 3278 14642 3330
rect 25678 3278 25730 3330
rect 28478 3278 28530 3330
rect 29710 3278 29762 3330
rect 65550 3278 65602 3330
rect 98142 3278 98194 3330
rect 122446 3278 122498 3330
rect 123342 3278 123394 3330
rect 124238 3278 124290 3330
rect 125134 3278 125186 3330
rect 126030 3278 126082 3330
rect 127598 3278 127650 3330
rect 128158 3278 128210 3330
rect 129390 3278 129442 3330
rect 130062 3278 130114 3330
rect 131182 3278 131234 3330
rect 132414 3278 132466 3330
rect 132974 3278 133026 3330
rect 133870 3278 133922 3330
rect 135998 3278 136050 3330
rect 136894 3278 136946 3330
rect 137790 3278 137842 3330
rect 139358 3278 139410 3330
rect 139918 3278 139970 3330
rect 140814 3278 140866 3330
rect 141710 3278 141762 3330
rect 142942 3278 142994 3330
rect 143838 3278 143890 3330
rect 144734 3278 144786 3330
rect 146862 3278 146914 3330
rect 147758 3278 147810 3330
rect 149550 3278 149602 3330
rect 150782 3278 150834 3330
rect 151678 3278 151730 3330
rect 152574 3278 152626 3330
rect 153470 3278 153522 3330
rect 154702 3278 154754 3330
rect 155598 3278 155650 3330
rect 156494 3278 156546 3330
rect 158622 3278 158674 3330
rect 159518 3278 159570 3330
rect 160414 3278 160466 3330
rect 161310 3278 161362 3330
rect 162542 3278 162594 3330
rect 163438 3278 163490 3330
rect 164334 3278 164386 3330
rect 165230 3278 165282 3330
rect 166462 3278 166514 3330
rect 167358 3278 167410 3330
rect 168254 3278 168306 3330
rect 169150 3278 169202 3330
rect 170382 3278 170434 3330
rect 171278 3278 171330 3330
rect 172174 3278 172226 3330
rect 173070 3278 173122 3330
rect 174302 3278 174354 3330
rect 174974 3278 175026 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 81278 3110 81330 3162
rect 81382 3110 81434 3162
rect 81486 3110 81538 3162
rect 111998 3110 112050 3162
rect 112102 3110 112154 3162
rect 112206 3110 112258 3162
rect 142718 3110 142770 3162
rect 142822 3110 142874 3162
rect 142926 3110 142978 3162
rect 173438 3110 173490 3162
rect 173542 3110 173594 3162
rect 173646 3110 173698 3162
rect 128718 2942 128770 2994
rect 129390 2942 129442 2994
rect 173406 1710 173458 1762
rect 174302 1710 174354 1762
<< metal2 >>
rect 1344 119200 1456 120000
rect 2912 119200 3024 120000
rect 4480 119200 4592 120000
rect 6048 119200 6160 120000
rect 7616 119200 7728 120000
rect 9184 119200 9296 120000
rect 10752 119200 10864 120000
rect 12320 119200 12432 120000
rect 13888 119200 14000 120000
rect 15456 119200 15568 120000
rect 17024 119200 17136 120000
rect 18592 119200 18704 120000
rect 20160 119200 20272 120000
rect 21728 119200 21840 120000
rect 23296 119200 23408 120000
rect 24864 119200 24976 120000
rect 26432 119200 26544 120000
rect 28000 119200 28112 120000
rect 29568 119200 29680 120000
rect 31136 119200 31248 120000
rect 32704 119200 32816 120000
rect 34272 119200 34384 120000
rect 35840 119200 35952 120000
rect 37408 119200 37520 120000
rect 38976 119200 39088 120000
rect 40544 119200 40656 120000
rect 42112 119200 42224 120000
rect 43680 119200 43792 120000
rect 45248 119200 45360 120000
rect 46816 119200 46928 120000
rect 48384 119200 48496 120000
rect 49952 119200 50064 120000
rect 51520 119200 51632 120000
rect 53088 119200 53200 120000
rect 54656 119200 54768 120000
rect 56224 119200 56336 120000
rect 57792 119200 57904 120000
rect 59360 119200 59472 120000
rect 60928 119200 61040 120000
rect 62496 119200 62608 120000
rect 64064 119200 64176 120000
rect 65632 119200 65744 120000
rect 67200 119200 67312 120000
rect 68768 119200 68880 120000
rect 70336 119200 70448 120000
rect 71904 119200 72016 120000
rect 73472 119200 73584 120000
rect 75040 119200 75152 120000
rect 76608 119200 76720 120000
rect 78176 119200 78288 120000
rect 79744 119200 79856 120000
rect 81312 119200 81424 120000
rect 82880 119200 82992 120000
rect 84448 119200 84560 120000
rect 86016 119200 86128 120000
rect 87584 119200 87696 120000
rect 89152 119200 89264 120000
rect 90720 119200 90832 120000
rect 92288 119200 92400 120000
rect 93856 119200 93968 120000
rect 95424 119200 95536 120000
rect 96992 119200 97104 120000
rect 98560 119200 98672 120000
rect 100128 119200 100240 120000
rect 101696 119200 101808 120000
rect 103264 119200 103376 120000
rect 104832 119200 104944 120000
rect 106400 119200 106512 120000
rect 107968 119200 108080 120000
rect 109536 119200 109648 120000
rect 111104 119200 111216 120000
rect 112672 119200 112784 120000
rect 114240 119200 114352 120000
rect 115808 119200 115920 120000
rect 117376 119200 117488 120000
rect 118944 119200 119056 120000
rect 120512 119200 120624 120000
rect 122080 119200 122192 120000
rect 123648 119200 123760 120000
rect 125216 119200 125328 120000
rect 126784 119200 126896 120000
rect 128352 119200 128464 120000
rect 129920 119200 130032 120000
rect 131488 119200 131600 120000
rect 133056 119200 133168 120000
rect 134624 119200 134736 120000
rect 136192 119200 136304 120000
rect 137760 119200 137872 120000
rect 139328 119200 139440 120000
rect 140896 119200 141008 120000
rect 142464 119200 142576 120000
rect 144032 119200 144144 120000
rect 145600 119200 145712 120000
rect 147168 119200 147280 120000
rect 148736 119200 148848 120000
rect 150304 119200 150416 120000
rect 151872 119200 151984 120000
rect 153440 119200 153552 120000
rect 155008 119200 155120 120000
rect 156576 119200 156688 120000
rect 158144 119200 158256 120000
rect 159712 119200 159824 120000
rect 161280 119200 161392 120000
rect 162848 119200 162960 120000
rect 164416 119200 164528 120000
rect 165984 119200 166096 120000
rect 167552 119200 167664 120000
rect 169120 119200 169232 120000
rect 170688 119200 170800 120000
rect 172256 119200 172368 120000
rect 173824 119200 173936 120000
rect 175392 119200 175504 120000
rect 176960 119200 177072 120000
rect 178528 119200 178640 120000
rect 2940 116564 2996 119200
rect 4508 117012 4564 119200
rect 4508 116946 4564 116956
rect 5964 117012 6020 117022
rect 4476 116844 4740 116854
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4476 116778 4740 116788
rect 2940 116498 2996 116508
rect 3388 116564 3444 116574
rect 3388 116470 3444 116508
rect 5964 116562 6020 116956
rect 7644 116676 7700 119200
rect 7644 116610 7700 116620
rect 8428 116676 8484 116686
rect 5964 116510 5966 116562
rect 6018 116510 6020 116562
rect 5964 116498 6020 116510
rect 8428 116562 8484 116620
rect 8428 116510 8430 116562
rect 8482 116510 8484 116562
rect 8428 116498 8484 116510
rect 9212 116564 9268 119200
rect 9212 116498 9268 116508
rect 10108 116564 10164 116574
rect 10108 116470 10164 116508
rect 4396 116450 4452 116462
rect 4396 116398 4398 116450
rect 4450 116398 4452 116450
rect 4396 115890 4452 116398
rect 4396 115838 4398 115890
rect 4450 115838 4452 115890
rect 4396 115826 4452 115838
rect 6748 116450 6804 116462
rect 6748 116398 6750 116450
rect 6802 116398 6804 116450
rect 4732 115668 4788 115678
rect 5180 115668 5236 115678
rect 4732 115666 5180 115668
rect 4732 115614 4734 115666
rect 4786 115614 5180 115666
rect 4732 115612 5180 115614
rect 4732 115602 4788 115612
rect 5180 115536 5236 115612
rect 6636 115556 6692 115566
rect 6748 115556 6804 116398
rect 7644 116450 7700 116462
rect 7644 116398 7646 116450
rect 7698 116398 7700 116450
rect 7532 115892 7588 115902
rect 7644 115892 7700 116398
rect 10892 116450 10948 116462
rect 10892 116398 10894 116450
rect 10946 116398 10948 116450
rect 10892 116228 10948 116398
rect 10892 116162 10948 116172
rect 11340 116228 11396 116238
rect 11340 116134 11396 116172
rect 7532 115890 7700 115892
rect 7532 115838 7534 115890
rect 7586 115838 7700 115890
rect 7532 115836 7700 115838
rect 12348 115892 12404 119200
rect 13916 117908 13972 119200
rect 13916 117852 14420 117908
rect 14364 116562 14420 117852
rect 14364 116510 14366 116562
rect 14418 116510 14420 116562
rect 14364 116498 14420 116510
rect 15372 116452 15428 116462
rect 15372 116450 15876 116452
rect 15372 116398 15374 116450
rect 15426 116398 15876 116450
rect 15372 116396 15876 116398
rect 15372 116386 15428 116396
rect 7532 115826 7588 115836
rect 12348 115826 12404 115836
rect 12684 116228 12740 116238
rect 12012 115778 12068 115790
rect 12012 115726 12014 115778
rect 12066 115726 12068 115778
rect 7196 115668 7252 115678
rect 7196 115574 7252 115612
rect 7980 115668 8036 115678
rect 6636 115554 6804 115556
rect 6636 115502 6638 115554
rect 6690 115502 6804 115554
rect 6636 115500 6804 115502
rect 4476 115276 4740 115286
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4476 115210 4740 115220
rect 4476 113708 4740 113718
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4476 113642 4740 113652
rect 4476 112140 4740 112150
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4476 112074 4740 112084
rect 4476 110572 4740 110582
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4476 110506 4740 110516
rect 4476 109004 4740 109014
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4476 108938 4740 108948
rect 6636 108388 6692 115500
rect 7980 114268 8036 115612
rect 11116 115668 11172 115678
rect 11116 115574 11172 115612
rect 11676 115668 11732 115678
rect 12012 115668 12068 115726
rect 12572 115668 12628 115678
rect 12012 115666 12628 115668
rect 12012 115614 12574 115666
rect 12626 115614 12628 115666
rect 12012 115612 12628 115614
rect 11676 115574 11732 115612
rect 12572 115602 12628 115612
rect 7980 114212 8148 114268
rect 6636 108322 6692 108332
rect 4476 107436 4740 107446
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4476 107370 4740 107380
rect 4476 105868 4740 105878
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4476 105802 4740 105812
rect 4476 104300 4740 104310
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4476 104234 4740 104244
rect 4476 102732 4740 102742
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4476 102666 4740 102676
rect 4476 101164 4740 101174
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4476 101098 4740 101108
rect 4476 99596 4740 99606
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4476 99530 4740 99540
rect 4476 98028 4740 98038
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4476 97962 4740 97972
rect 4476 96460 4740 96470
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4476 96394 4740 96404
rect 4476 94892 4740 94902
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4476 94826 4740 94836
rect 4476 93324 4740 93334
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4476 93258 4740 93268
rect 4476 91756 4740 91766
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4476 91690 4740 91700
rect 4476 90188 4740 90198
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4476 90122 4740 90132
rect 4476 88620 4740 88630
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4476 88554 4740 88564
rect 4476 87052 4740 87062
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4476 86986 4740 86996
rect 4476 85484 4740 85494
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4476 85418 4740 85428
rect 4476 83916 4740 83926
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4476 83850 4740 83860
rect 4476 82348 4740 82358
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4476 82282 4740 82292
rect 4476 80780 4740 80790
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4476 80714 4740 80724
rect 4476 79212 4740 79222
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4476 79146 4740 79156
rect 4476 77644 4740 77654
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4476 77578 4740 77588
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 8092 20188 8148 114212
rect 12684 102508 12740 116172
rect 15820 116226 15876 116396
rect 15820 116174 15822 116226
rect 15874 116174 15876 116226
rect 13244 115892 13300 115902
rect 13244 115554 13300 115836
rect 13244 115502 13246 115554
rect 13298 115502 13300 115554
rect 13244 115490 13300 115502
rect 12572 102452 12740 102508
rect 8988 20244 9044 20254
rect 8092 20132 8372 20188
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5964 8484 6020 8494
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 5852 3444 5908 3454
rect 5852 3350 5908 3388
rect 5964 800 6020 8428
rect 8204 5908 8260 5918
rect 7980 5796 8036 5806
rect 8204 5796 8260 5852
rect 7980 5794 8260 5796
rect 7980 5742 7982 5794
rect 8034 5742 8260 5794
rect 7980 5740 8260 5742
rect 7980 5730 8036 5740
rect 7644 5122 7700 5134
rect 7644 5070 7646 5122
rect 7698 5070 7700 5122
rect 7084 4900 7140 4910
rect 7644 4900 7700 5070
rect 7868 5124 7924 5134
rect 7868 5010 7924 5068
rect 7868 4958 7870 5010
rect 7922 4958 7924 5010
rect 7868 4946 7924 4958
rect 7084 4898 7700 4900
rect 7084 4846 7086 4898
rect 7138 4846 7700 4898
rect 7084 4844 7700 4846
rect 7084 4834 7140 4844
rect 6860 4226 6916 4238
rect 7532 4228 7588 4238
rect 6860 4174 6862 4226
rect 6914 4174 6916 4226
rect 6860 4116 6916 4174
rect 6860 4050 6916 4060
rect 7084 4226 7588 4228
rect 7084 4174 7534 4226
rect 7586 4174 7588 4226
rect 7084 4172 7588 4174
rect 6524 3554 6580 3566
rect 6524 3502 6526 3554
rect 6578 3502 6580 3554
rect 6524 3444 6580 3502
rect 6524 800 6580 3388
rect 7084 800 7140 4172
rect 7532 4162 7588 4172
rect 7644 800 7700 4844
rect 8204 800 8260 5740
rect 8316 3666 8372 20132
rect 8428 6018 8484 6030
rect 8428 5966 8430 6018
rect 8482 5966 8484 6018
rect 8428 5234 8484 5966
rect 8652 5908 8708 5918
rect 8652 5814 8708 5852
rect 8988 5346 9044 20188
rect 12572 19348 12628 102452
rect 12572 19282 12628 19292
rect 15148 16884 15204 16894
rect 14924 7362 14980 7374
rect 14924 7310 14926 7362
rect 14978 7310 14980 7362
rect 14924 6692 14980 7310
rect 14700 6636 14980 6692
rect 14588 6578 14644 6590
rect 14588 6526 14590 6578
rect 14642 6526 14644 6578
rect 14140 6468 14196 6478
rect 14588 6468 14644 6526
rect 14140 6466 14644 6468
rect 14140 6414 14142 6466
rect 14194 6414 14644 6466
rect 14140 6412 14644 6414
rect 11564 6132 11620 6142
rect 9660 5796 9716 5806
rect 8988 5294 8990 5346
rect 9042 5294 9044 5346
rect 8988 5282 9044 5294
rect 9548 5794 9716 5796
rect 9548 5742 9662 5794
rect 9714 5742 9716 5794
rect 9548 5740 9716 5742
rect 8428 5182 8430 5234
rect 8482 5182 8484 5234
rect 8428 5170 8484 5182
rect 8652 5124 8708 5134
rect 8652 5030 8708 5068
rect 9548 5010 9604 5740
rect 9660 5730 9716 5740
rect 11228 5794 11284 5806
rect 11228 5742 11230 5794
rect 11282 5742 11284 5794
rect 10668 5572 10724 5582
rect 9548 4958 9550 5010
rect 9602 4958 9604 5010
rect 8540 4338 8596 4350
rect 8540 4286 8542 4338
rect 8594 4286 8596 4338
rect 8540 4116 8596 4286
rect 9100 4228 9156 4238
rect 9100 4134 9156 4172
rect 8540 4050 8596 4060
rect 8316 3614 8318 3666
rect 8370 3614 8372 3666
rect 8316 980 8372 3614
rect 9548 3556 9604 4958
rect 9884 5012 9940 5022
rect 9884 4918 9940 4956
rect 10444 4564 10500 4574
rect 10444 4470 10500 4508
rect 10108 4340 10164 4350
rect 8316 914 8372 924
rect 8764 3500 9604 3556
rect 9884 4338 10164 4340
rect 9884 4286 10110 4338
rect 10162 4286 10164 4338
rect 9884 4284 10164 4286
rect 9884 4228 9940 4284
rect 10108 4274 10164 4284
rect 8764 800 8820 3500
rect 9884 800 9940 4172
rect 10332 3668 10388 3678
rect 10332 3666 10500 3668
rect 10332 3614 10334 3666
rect 10386 3614 10500 3666
rect 10332 3612 10500 3614
rect 10332 3602 10388 3612
rect 10444 800 10500 3612
rect 10668 3556 10724 5516
rect 11228 5572 11284 5742
rect 11228 5506 11284 5516
rect 11228 5010 11284 5022
rect 11228 4958 11230 5010
rect 11282 4958 11284 5010
rect 10780 4898 10836 4910
rect 10780 4846 10782 4898
rect 10834 4846 10836 4898
rect 10780 4564 10836 4846
rect 11228 4564 11284 4958
rect 11564 5010 11620 6076
rect 13468 6020 13524 6030
rect 13468 5926 13524 5964
rect 13244 5906 13300 5918
rect 13244 5854 13246 5906
rect 13298 5854 13300 5906
rect 11788 5794 11844 5806
rect 11788 5742 11790 5794
rect 11842 5742 11844 5794
rect 11564 4958 11566 5010
rect 11618 4958 11620 5010
rect 11564 4946 11620 4958
rect 11676 5124 11732 5134
rect 10780 4508 11284 4564
rect 10780 3556 10836 3566
rect 10668 3554 10836 3556
rect 10668 3502 10782 3554
rect 10834 3502 10836 3554
rect 10668 3500 10836 3502
rect 10780 3490 10836 3500
rect 11004 800 11060 4508
rect 11452 4450 11508 4462
rect 11452 4398 11454 4450
rect 11506 4398 11508 4450
rect 11228 4338 11284 4350
rect 11228 4286 11230 4338
rect 11282 4286 11284 4338
rect 11228 3444 11284 4286
rect 11452 3780 11508 4398
rect 11452 3714 11508 3724
rect 11228 3378 11284 3388
rect 11676 3554 11732 5068
rect 11676 3502 11678 3554
rect 11730 3502 11732 3554
rect 11676 2660 11732 3502
rect 11788 3444 11844 5742
rect 12684 5796 12740 5806
rect 13244 5796 13300 5854
rect 12684 5794 13300 5796
rect 12684 5742 12686 5794
rect 12738 5742 13300 5794
rect 12684 5740 13300 5742
rect 12684 5730 12740 5740
rect 12012 5124 12068 5134
rect 12012 5030 12068 5068
rect 12908 5124 12964 5134
rect 12908 5010 12964 5068
rect 12908 4958 12910 5010
rect 12962 4958 12964 5010
rect 12908 4946 12964 4958
rect 12572 4900 12628 4910
rect 12572 4898 12852 4900
rect 12572 4846 12574 4898
rect 12626 4846 12852 4898
rect 12572 4844 12852 4846
rect 12572 4834 12628 4844
rect 12796 4450 12852 4844
rect 12796 4398 12798 4450
rect 12850 4398 12852 4450
rect 12796 4386 12852 4398
rect 12124 4338 12180 4350
rect 12124 4286 12126 4338
rect 12178 4286 12180 4338
rect 12124 3668 12180 4286
rect 12124 3602 12180 3612
rect 12572 3668 12628 3678
rect 12572 3666 12740 3668
rect 12572 3614 12574 3666
rect 12626 3614 12740 3666
rect 12572 3612 12740 3614
rect 12572 3602 12628 3612
rect 11788 3378 11844 3388
rect 12124 3444 12180 3454
rect 11676 2594 11732 2604
rect 12124 800 12180 3388
rect 12684 800 12740 3612
rect 13244 800 13300 5740
rect 14028 5906 14084 5918
rect 14028 5854 14030 5906
rect 14082 5854 14084 5906
rect 13692 5236 13748 5246
rect 13692 5142 13748 5180
rect 14028 5012 14084 5854
rect 14028 4946 14084 4956
rect 14140 4340 14196 6412
rect 14364 6018 14420 6030
rect 14364 5966 14366 6018
rect 14418 5966 14420 6018
rect 14364 5908 14420 5966
rect 14364 5842 14420 5852
rect 14588 5348 14644 5358
rect 14588 5254 14644 5292
rect 14252 5124 14308 5134
rect 14252 5030 14308 5068
rect 14140 4284 14420 4340
rect 13804 3668 13860 3678
rect 13804 3574 13860 3612
rect 14252 3556 14308 3566
rect 14252 3462 14308 3500
rect 14364 800 14420 4284
rect 14700 3556 14756 6636
rect 14924 6468 14980 6478
rect 14924 6374 14980 6412
rect 14812 6244 14868 6254
rect 14812 5236 14868 6188
rect 15148 6132 15204 16828
rect 15820 8708 15876 116174
rect 17052 115892 17108 119200
rect 18620 117908 18676 119200
rect 18620 117852 19124 117908
rect 19068 116562 19124 117852
rect 21756 117572 21812 119200
rect 21756 117516 22260 117572
rect 19068 116510 19070 116562
rect 19122 116510 19124 116562
rect 19068 116498 19124 116510
rect 22204 116562 22260 117516
rect 22204 116510 22206 116562
rect 22258 116510 22260 116562
rect 22204 116498 22260 116510
rect 23324 116564 23380 119200
rect 26460 117236 26516 119200
rect 26460 117170 26516 117180
rect 27356 117236 27412 117246
rect 23548 116564 23604 116574
rect 23324 116562 23604 116564
rect 23324 116510 23550 116562
rect 23602 116510 23604 116562
rect 23324 116508 23604 116510
rect 23548 116498 23604 116508
rect 27356 116562 27412 117180
rect 27356 116510 27358 116562
rect 27410 116510 27412 116562
rect 27356 116498 27412 116510
rect 28028 116564 28084 119200
rect 30492 117010 30548 117022
rect 30492 116958 30494 117010
rect 30546 116958 30548 117010
rect 28028 116498 28084 116508
rect 29484 116564 29540 116574
rect 29484 116470 29540 116508
rect 17052 115826 17108 115836
rect 18060 116452 18116 116462
rect 16940 115778 16996 115790
rect 16940 115726 16942 115778
rect 16994 115726 16996 115778
rect 16044 115668 16100 115678
rect 16044 115574 16100 115612
rect 16716 115668 16772 115678
rect 16940 115668 16996 115726
rect 17724 115668 17780 115678
rect 16940 115666 17780 115668
rect 16940 115614 17726 115666
rect 17778 115614 17780 115666
rect 16940 115612 17780 115614
rect 16716 115574 16772 115612
rect 17724 115602 17780 115612
rect 18060 20188 18116 116396
rect 19852 116452 19908 116462
rect 19852 116358 19908 116396
rect 20524 116452 20580 116462
rect 20524 116358 20580 116396
rect 21756 116450 21812 116462
rect 21756 116398 21758 116450
rect 21810 116398 21812 116450
rect 19836 116060 20100 116070
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 19836 115994 20100 116004
rect 18620 115892 18676 115902
rect 18620 115778 18676 115836
rect 21756 115890 21812 116398
rect 24556 116452 24612 116462
rect 26684 116452 26740 116462
rect 24556 116450 24836 116452
rect 24556 116398 24558 116450
rect 24610 116398 24836 116450
rect 24556 116396 24836 116398
rect 24556 116386 24612 116396
rect 21756 115838 21758 115890
rect 21810 115838 21812 115890
rect 21756 115826 21812 115838
rect 24780 116228 24836 116396
rect 26460 116450 26740 116452
rect 26460 116398 26686 116450
rect 26738 116398 26740 116450
rect 26460 116396 26740 116398
rect 25228 116228 25284 116238
rect 24780 116226 25284 116228
rect 24780 116174 25230 116226
rect 25282 116174 25284 116226
rect 24780 116172 25284 116174
rect 18620 115726 18622 115778
rect 18674 115726 18676 115778
rect 18620 115714 18676 115726
rect 20860 115668 20916 115678
rect 20860 115574 20916 115612
rect 21532 115668 21588 115678
rect 21532 115574 21588 115612
rect 19836 114492 20100 114502
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 19836 114426 20100 114436
rect 19836 112924 20100 112934
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 19836 112858 20100 112868
rect 19836 111356 20100 111366
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 19836 111290 20100 111300
rect 19836 109788 20100 109798
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 19836 109722 20100 109732
rect 19836 108220 20100 108230
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 19836 108154 20100 108164
rect 19836 106652 20100 106662
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 19836 106586 20100 106596
rect 19836 105084 20100 105094
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 19836 105018 20100 105028
rect 19836 103516 20100 103526
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 19836 103450 20100 103460
rect 19836 101948 20100 101958
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 19836 101882 20100 101892
rect 19836 100380 20100 100390
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 19836 100314 20100 100324
rect 19836 98812 20100 98822
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 19836 98746 20100 98756
rect 19836 97244 20100 97254
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 19836 97178 20100 97188
rect 19836 95676 20100 95686
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 19836 95610 20100 95620
rect 19836 94108 20100 94118
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 19836 94042 20100 94052
rect 19836 92540 20100 92550
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 19836 92474 20100 92484
rect 19836 90972 20100 90982
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 19836 90906 20100 90916
rect 19836 89404 20100 89414
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 19836 89338 20100 89348
rect 19836 87836 20100 87846
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 19836 87770 20100 87780
rect 19836 86268 20100 86278
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 19836 86202 20100 86212
rect 19836 84700 20100 84710
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 19836 84634 20100 84644
rect 19836 83132 20100 83142
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 19836 83066 20100 83076
rect 19836 81564 20100 81574
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 19836 81498 20100 81508
rect 19836 79996 20100 80006
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 19836 79930 20100 79940
rect 19836 78428 20100 78438
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 19836 78362 20100 78372
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 18060 20132 18228 20188
rect 15484 6466 15540 6478
rect 15484 6414 15486 6466
rect 15538 6414 15540 6466
rect 15260 6132 15316 6142
rect 15148 6130 15316 6132
rect 15148 6078 15262 6130
rect 15314 6078 15316 6130
rect 15148 6076 15316 6078
rect 15260 6066 15316 6076
rect 14924 6020 14980 6030
rect 14924 5926 14980 5964
rect 15036 6018 15092 6030
rect 15036 5966 15038 6018
rect 15090 5966 15092 6018
rect 14812 5010 14868 5180
rect 15036 5236 15092 5966
rect 15036 5170 15092 5180
rect 15484 5908 15540 6414
rect 15820 6466 15876 8652
rect 16828 18564 16884 18574
rect 16380 7362 16436 7374
rect 16380 7310 16382 7362
rect 16434 7310 16436 7362
rect 16380 7252 16436 7310
rect 15820 6414 15822 6466
rect 15874 6414 15876 6466
rect 15708 5908 15764 5918
rect 15484 5906 15764 5908
rect 15484 5854 15710 5906
rect 15762 5854 15764 5906
rect 15484 5852 15764 5854
rect 15148 5012 15204 5022
rect 14812 4958 14814 5010
rect 14866 4958 14868 5010
rect 14812 4946 14868 4958
rect 14924 5010 15204 5012
rect 14924 4958 15150 5010
rect 15202 4958 15204 5010
rect 14924 4956 15204 4958
rect 14924 4226 14980 4956
rect 15148 4946 15204 4956
rect 14924 4174 14926 4226
rect 14978 4174 14980 4226
rect 14924 3556 14980 4174
rect 15148 3556 15204 3566
rect 14924 3554 15204 3556
rect 14924 3502 15150 3554
rect 15202 3502 15204 3554
rect 14924 3500 15204 3502
rect 14700 3490 14756 3500
rect 15148 3490 15204 3500
rect 14812 3444 14868 3454
rect 14868 3388 14980 3444
rect 14812 3378 14868 3388
rect 14588 3332 14644 3342
rect 14588 3238 14644 3276
rect 14924 800 14980 3388
rect 15484 800 15540 5852
rect 15708 5842 15764 5852
rect 15820 5348 15876 6414
rect 15820 5282 15876 5292
rect 15932 7196 16436 7252
rect 15820 4340 15876 4350
rect 15932 4340 15988 7196
rect 16380 6466 16436 6478
rect 16380 6414 16382 6466
rect 16434 6414 16436 6466
rect 16380 6356 16436 6414
rect 16380 6290 16436 6300
rect 16044 6132 16100 6142
rect 16716 6132 16772 6142
rect 16044 6130 16772 6132
rect 16044 6078 16046 6130
rect 16098 6078 16718 6130
rect 16770 6078 16772 6130
rect 16044 6076 16772 6078
rect 16828 6132 16884 18508
rect 16940 6468 16996 6478
rect 16940 6466 17220 6468
rect 16940 6414 16942 6466
rect 16994 6414 17220 6466
rect 16940 6412 17220 6414
rect 16940 6402 16996 6412
rect 16940 6132 16996 6142
rect 16828 6130 16996 6132
rect 16828 6078 16942 6130
rect 16994 6078 16996 6130
rect 16828 6076 16996 6078
rect 16044 6066 16100 6076
rect 16716 6066 16772 6076
rect 16940 6066 16996 6076
rect 16604 5908 16660 5918
rect 16604 5814 16660 5852
rect 16044 5348 16100 5358
rect 16044 4562 16100 5292
rect 16044 4510 16046 4562
rect 16098 4510 16100 4562
rect 16044 4498 16100 4510
rect 16156 5122 16212 5134
rect 16828 5124 16884 5134
rect 16156 5070 16158 5122
rect 16210 5070 16212 5122
rect 15820 4338 15988 4340
rect 15820 4286 15822 4338
rect 15874 4286 15988 4338
rect 15820 4284 15988 4286
rect 15820 4004 15876 4284
rect 16156 4228 16212 5070
rect 16604 5122 16884 5124
rect 16604 5070 16830 5122
rect 16882 5070 16884 5122
rect 16604 5068 16884 5070
rect 16604 4562 16660 5068
rect 16828 5058 16884 5068
rect 16604 4510 16606 4562
rect 16658 4510 16660 4562
rect 16604 4498 16660 4510
rect 17164 4452 17220 6412
rect 17388 6466 17444 6478
rect 17388 6414 17390 6466
rect 17442 6414 17444 6466
rect 17388 6356 17444 6414
rect 17388 5908 17444 6300
rect 17724 6466 17780 6478
rect 17724 6414 17726 6466
rect 17778 6414 17780 6466
rect 17724 6244 17780 6414
rect 17724 6178 17780 6188
rect 18172 6466 18228 20132
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 23100 18676 23156 18686
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 21980 13636 22036 13646
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 18620 10164 18676 10174
rect 18284 7474 18340 7486
rect 18284 7422 18286 7474
rect 18338 7422 18340 7474
rect 18284 7364 18340 7422
rect 18284 7298 18340 7308
rect 18172 6414 18174 6466
rect 18226 6414 18228 6466
rect 17388 5842 17444 5852
rect 17836 5684 17892 5694
rect 17164 4386 17220 4396
rect 17388 5682 17892 5684
rect 17388 5630 17838 5682
rect 17890 5630 17892 5682
rect 17388 5628 17892 5630
rect 16940 4338 16996 4350
rect 16940 4286 16942 4338
rect 16994 4286 16996 4338
rect 16940 4228 16996 4286
rect 17388 4228 17444 5628
rect 17836 5618 17892 5628
rect 18172 5682 18228 6414
rect 18396 6244 18452 6254
rect 18396 6020 18452 6188
rect 18396 5888 18452 5964
rect 18172 5630 18174 5682
rect 18226 5630 18228 5682
rect 16940 4172 17444 4228
rect 17836 4228 17892 4238
rect 16156 4162 16212 4172
rect 17836 4134 17892 4172
rect 15820 3938 15876 3948
rect 17724 4004 17780 4014
rect 16604 3556 16660 3566
rect 16044 3444 16100 3454
rect 16044 3350 16100 3388
rect 16604 800 16660 3500
rect 17164 3444 17220 3454
rect 17164 800 17220 3388
rect 17724 800 17780 3948
rect 17836 3444 17892 3454
rect 17836 3350 17892 3388
rect 18172 2772 18228 5630
rect 18620 4564 18676 10108
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 8146 19684 8158
rect 19628 8094 19630 8146
rect 19682 8094 19684 8146
rect 19292 8036 19348 8046
rect 18956 8034 19348 8036
rect 18956 7982 19294 8034
rect 19346 7982 19348 8034
rect 18956 7980 19348 7982
rect 18956 7586 19012 7980
rect 19292 7970 19348 7980
rect 18956 7534 18958 7586
rect 19010 7534 19012 7586
rect 18956 7522 19012 7534
rect 19292 7364 19348 7374
rect 18732 6578 18788 6590
rect 18732 6526 18734 6578
rect 18786 6526 18788 6578
rect 18732 5348 18788 6526
rect 18844 6466 18900 6478
rect 18844 6414 18846 6466
rect 18898 6414 18900 6466
rect 18844 6356 18900 6414
rect 18844 6290 18900 6300
rect 19068 6466 19124 6478
rect 19068 6414 19070 6466
rect 19122 6414 19124 6466
rect 18732 5282 18788 5292
rect 18956 6018 19012 6030
rect 18956 5966 18958 6018
rect 19010 5966 19012 6018
rect 18956 5234 19012 5966
rect 18956 5182 18958 5234
rect 19010 5182 19012 5234
rect 18732 4564 18788 4574
rect 18620 4562 18788 4564
rect 18620 4510 18734 4562
rect 18786 4510 18788 4562
rect 18620 4508 18788 4510
rect 18732 4498 18788 4508
rect 18396 4452 18452 4462
rect 18396 4340 18452 4396
rect 18396 4338 18564 4340
rect 18396 4286 18398 4338
rect 18450 4286 18564 4338
rect 18396 4284 18564 4286
rect 18396 4274 18452 4284
rect 18508 3332 18564 4284
rect 18732 3556 18788 3566
rect 18956 3556 19012 5182
rect 19068 5236 19124 6414
rect 19068 5170 19124 5180
rect 19180 6356 19236 6366
rect 19180 4900 19236 6300
rect 19180 4834 19236 4844
rect 19292 4338 19348 7308
rect 19628 6914 19684 8094
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 21084 7362 21140 7374
rect 21084 7310 21086 7362
rect 21138 7310 21140 7362
rect 19628 6862 19630 6914
rect 19682 6862 19684 6914
rect 19628 6850 19684 6862
rect 19964 6916 20020 6926
rect 19964 6822 20020 6860
rect 20636 6690 20692 6702
rect 20636 6638 20638 6690
rect 20690 6638 20692 6690
rect 20188 6580 20244 6590
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20188 6132 20244 6524
rect 20636 6580 20692 6638
rect 20636 6514 20692 6524
rect 20748 6580 20804 6590
rect 21084 6580 21140 7310
rect 21532 7364 21588 7374
rect 21532 7270 21588 7308
rect 21980 7362 22036 13580
rect 22764 9380 22820 9390
rect 21980 7310 21982 7362
rect 22034 7310 22036 7362
rect 21980 7252 22036 7310
rect 22428 7364 22484 7374
rect 22428 7270 22484 7308
rect 21980 6916 22036 7196
rect 21980 6850 22036 6860
rect 22092 7140 22148 7150
rect 20748 6578 21140 6580
rect 20748 6526 20750 6578
rect 20802 6526 21140 6578
rect 20748 6524 21140 6526
rect 21532 6580 21588 6590
rect 20076 6076 20244 6132
rect 20076 6020 20132 6076
rect 20300 6020 20356 6030
rect 20076 5954 20132 5964
rect 20188 6018 20356 6020
rect 20188 5966 20302 6018
rect 20354 5966 20356 6018
rect 20188 5964 20356 5966
rect 19852 5796 19908 5806
rect 19852 5702 19908 5740
rect 19852 5236 19908 5246
rect 19292 4286 19294 4338
rect 19346 4286 19348 4338
rect 19292 3668 19348 4286
rect 19292 3602 19348 3612
rect 19404 5234 19908 5236
rect 19404 5182 19854 5234
rect 19906 5182 19908 5234
rect 19404 5180 19908 5182
rect 18732 3554 19012 3556
rect 18732 3502 18734 3554
rect 18786 3502 19012 3554
rect 18732 3500 19012 3502
rect 18732 3490 18788 3500
rect 18508 3276 18900 3332
rect 18172 2706 18228 2716
rect 18844 800 18900 3276
rect 19404 800 19460 5180
rect 19852 5170 19908 5180
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20188 4564 20244 5964
rect 20300 5954 20356 5964
rect 20636 5906 20692 5918
rect 20636 5854 20638 5906
rect 20690 5854 20692 5906
rect 20076 4508 20244 4564
rect 20524 5796 20580 5806
rect 20076 4450 20132 4508
rect 20076 4398 20078 4450
rect 20130 4398 20132 4450
rect 20076 4386 20132 4398
rect 19740 3444 19796 3454
rect 19740 3350 19796 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20524 800 20580 5740
rect 20636 4676 20692 5854
rect 20748 5122 20804 6524
rect 21532 6486 21588 6524
rect 21532 6020 21588 6030
rect 21532 6018 21812 6020
rect 21532 5966 21534 6018
rect 21586 5966 21812 6018
rect 21532 5964 21812 5966
rect 21532 5954 21588 5964
rect 21196 5906 21252 5918
rect 21196 5854 21198 5906
rect 21250 5854 21252 5906
rect 21196 5796 21252 5854
rect 21196 5730 21252 5740
rect 20748 5070 20750 5122
rect 20802 5070 20804 5122
rect 20748 5058 20804 5070
rect 21644 5236 21700 5246
rect 20636 4620 21588 4676
rect 21532 3778 21588 4620
rect 21532 3726 21534 3778
rect 21586 3726 21588 3778
rect 21532 3714 21588 3726
rect 20636 3556 20692 3566
rect 20636 3462 20692 3500
rect 21084 3444 21140 3454
rect 21084 800 21140 3388
rect 21644 1652 21700 5180
rect 21644 1586 21700 1596
rect 21756 1204 21812 5964
rect 21868 5236 21924 5246
rect 21868 5142 21924 5180
rect 22092 5012 22148 7084
rect 22540 6580 22596 6590
rect 22652 6580 22708 6590
rect 22596 6578 22708 6580
rect 22596 6526 22654 6578
rect 22706 6526 22708 6578
rect 22596 6524 22708 6526
rect 22204 6466 22260 6478
rect 22204 6414 22206 6466
rect 22258 6414 22260 6466
rect 22204 5908 22260 6414
rect 22428 5908 22484 5918
rect 22204 5906 22484 5908
rect 22204 5854 22430 5906
rect 22482 5854 22484 5906
rect 22204 5852 22484 5854
rect 21868 4956 22148 5012
rect 21868 3778 21924 4956
rect 22204 4226 22260 4238
rect 22204 4174 22206 4226
rect 22258 4174 22260 4226
rect 22204 4116 22260 4174
rect 21868 3726 21870 3778
rect 21922 3726 21924 3778
rect 21868 3714 21924 3726
rect 21980 4060 22260 4116
rect 21980 3556 22036 4060
rect 22428 4004 22484 5852
rect 21980 3490 22036 3500
rect 22204 3948 22484 4004
rect 21756 1138 21812 1148
rect 22204 800 22260 3948
rect 22428 3556 22484 3566
rect 22428 3442 22484 3500
rect 22540 3554 22596 6524
rect 22652 6514 22708 6524
rect 22764 6130 22820 9324
rect 22876 7362 22932 7374
rect 22876 7310 22878 7362
rect 22930 7310 22932 7362
rect 22876 6580 22932 7310
rect 22876 6514 22932 6524
rect 22764 6078 22766 6130
rect 22818 6078 22820 6130
rect 22764 6066 22820 6078
rect 22540 3502 22542 3554
rect 22594 3502 22596 3554
rect 22540 3490 22596 3502
rect 22652 5010 22708 5022
rect 22652 4958 22654 5010
rect 22706 4958 22708 5010
rect 22428 3390 22430 3442
rect 22482 3390 22484 3442
rect 22428 3378 22484 3390
rect 22652 2548 22708 4958
rect 23100 4562 23156 18620
rect 24444 12852 24500 12862
rect 23436 7364 23492 7374
rect 23324 7362 23492 7364
rect 23324 7310 23438 7362
rect 23490 7310 23492 7362
rect 23324 7308 23492 7310
rect 23212 6466 23268 6478
rect 23212 6414 23214 6466
rect 23266 6414 23268 6466
rect 23212 6356 23268 6414
rect 23212 6290 23268 6300
rect 23100 4510 23102 4562
rect 23154 4510 23156 4562
rect 23100 4498 23156 4510
rect 22876 4340 22932 4350
rect 22876 4246 22932 4284
rect 23324 4340 23380 7308
rect 23436 7298 23492 7308
rect 23884 7362 23940 7374
rect 23884 7310 23886 7362
rect 23938 7310 23940 7362
rect 23548 6356 23604 6366
rect 23548 6130 23604 6300
rect 23548 6078 23550 6130
rect 23602 6078 23604 6130
rect 23548 6066 23604 6078
rect 23884 5908 23940 7310
rect 24220 7362 24276 7374
rect 24220 7310 24222 7362
rect 24274 7310 24276 7362
rect 24220 7140 24276 7310
rect 24220 7074 24276 7084
rect 24332 7252 24388 7262
rect 24108 6692 24164 6702
rect 24108 6690 24276 6692
rect 24108 6638 24110 6690
rect 24162 6638 24276 6690
rect 24108 6636 24276 6638
rect 24108 6626 24164 6636
rect 24108 5908 24164 5918
rect 23884 5906 24164 5908
rect 23884 5854 24110 5906
rect 24162 5854 24164 5906
rect 23884 5852 24164 5854
rect 24220 5908 24276 6636
rect 24332 6578 24388 7196
rect 24332 6526 24334 6578
rect 24386 6526 24388 6578
rect 24332 6514 24388 6526
rect 24444 6130 24500 12796
rect 24444 6078 24446 6130
rect 24498 6078 24500 6130
rect 24444 6066 24500 6078
rect 24780 6466 24836 116172
rect 25228 116162 25284 116172
rect 26460 115890 26516 116396
rect 26684 116386 26740 116396
rect 30492 116450 30548 116958
rect 31164 116676 31220 119200
rect 31164 116610 31220 116620
rect 31612 117010 31668 117022
rect 31612 116958 31614 117010
rect 31666 116958 31668 117010
rect 30492 116398 30494 116450
rect 30546 116398 30548 116450
rect 30492 116386 30548 116398
rect 31164 116450 31220 116462
rect 31164 116398 31166 116450
rect 31218 116398 31220 116450
rect 26460 115838 26462 115890
rect 26514 115838 26516 115890
rect 26460 115826 26516 115838
rect 31164 115890 31220 116398
rect 31164 115838 31166 115890
rect 31218 115838 31220 115890
rect 31164 115826 31220 115838
rect 31612 115890 31668 116958
rect 31948 116676 32004 116686
rect 31948 116562 32004 116620
rect 31948 116510 31950 116562
rect 32002 116510 32004 116562
rect 31948 116498 32004 116510
rect 32732 116564 32788 119200
rect 35196 116844 35460 116854
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35196 116778 35460 116788
rect 32732 116498 32788 116508
rect 33628 116564 33684 116574
rect 33628 116470 33684 116508
rect 34412 116452 34468 116462
rect 34412 116450 34916 116452
rect 34412 116398 34414 116450
rect 34466 116398 34916 116450
rect 34412 116396 34916 116398
rect 34412 116386 34468 116396
rect 31612 115838 31614 115890
rect 31666 115838 31668 115890
rect 25564 115668 25620 115678
rect 25564 115574 25620 115612
rect 26236 115668 26292 115678
rect 26236 115574 26292 115612
rect 30268 115668 30324 115678
rect 30268 115574 30324 115612
rect 30940 115668 30996 115678
rect 30940 115574 30996 115612
rect 25788 22596 25844 22606
rect 25788 8428 25844 22540
rect 31612 20188 31668 115838
rect 34860 116226 34916 116396
rect 34860 116174 34862 116226
rect 34914 116174 34916 116226
rect 34636 115668 34692 115678
rect 34636 115574 34692 115612
rect 31276 20132 31668 20188
rect 33628 22484 33684 22494
rect 25564 8372 25844 8428
rect 26908 16772 26964 16782
rect 24780 6414 24782 6466
rect 24834 6414 24836 6466
rect 24780 5908 24836 6414
rect 25340 6468 25396 6478
rect 25340 6466 25508 6468
rect 25340 6414 25342 6466
rect 25394 6414 25508 6466
rect 25340 6412 25508 6414
rect 25340 6402 25396 6412
rect 24892 6132 24948 6142
rect 24892 6038 24948 6076
rect 24220 5852 24836 5908
rect 23772 5236 23828 5246
rect 23436 5122 23492 5134
rect 23436 5070 23438 5122
rect 23490 5070 23492 5122
rect 23436 4452 23492 5070
rect 23436 4386 23492 4396
rect 23324 4274 23380 4284
rect 23772 4338 23828 5180
rect 23996 4452 24052 5852
rect 24108 5842 24164 5852
rect 23772 4286 23774 4338
rect 23826 4286 23828 4338
rect 23772 4274 23828 4286
rect 23884 4396 24052 4452
rect 24108 5234 24164 5246
rect 24108 5182 24110 5234
rect 24162 5182 24164 5234
rect 23660 3444 23716 3454
rect 23660 3350 23716 3388
rect 22652 2492 22820 2548
rect 22764 800 22820 2492
rect 23884 800 23940 4396
rect 24108 3556 24164 5182
rect 24108 3490 24164 3500
rect 24444 4226 24500 4238
rect 24444 4174 24446 4226
rect 24498 4174 24500 4226
rect 24444 800 24500 4174
rect 24556 3556 24612 3566
rect 24556 3462 24612 3500
rect 24780 1092 24836 5852
rect 25340 4340 25396 4350
rect 25340 3220 25396 4284
rect 25452 3780 25508 6412
rect 25452 3554 25508 3724
rect 25452 3502 25454 3554
rect 25506 3502 25508 3554
rect 25452 3490 25508 3502
rect 25564 3332 25620 8372
rect 26796 8036 26852 8046
rect 26460 8034 26852 8036
rect 26460 7982 26798 8034
rect 26850 7982 26852 8034
rect 26460 7980 26852 7982
rect 26460 7586 26516 7980
rect 26796 7970 26852 7980
rect 26460 7534 26462 7586
rect 26514 7534 26516 7586
rect 26460 7522 26516 7534
rect 26796 7812 26852 7822
rect 25676 7474 25732 7486
rect 25676 7422 25678 7474
rect 25730 7422 25732 7474
rect 25676 7364 25732 7422
rect 25676 6132 25732 7308
rect 25900 6692 25956 6702
rect 25900 6690 26740 6692
rect 25900 6638 25902 6690
rect 25954 6638 26740 6690
rect 25900 6636 26740 6638
rect 25900 6626 25956 6636
rect 26124 6468 26180 6478
rect 26124 6466 26516 6468
rect 26124 6414 26126 6466
rect 26178 6414 26516 6466
rect 26124 6412 26516 6414
rect 26124 6402 26180 6412
rect 25676 5906 25732 6076
rect 26460 6018 26516 6412
rect 26460 5966 26462 6018
rect 26514 5966 26516 6018
rect 26460 5954 26516 5966
rect 25676 5854 25678 5906
rect 25730 5854 25732 5906
rect 25676 5842 25732 5854
rect 26236 5012 26292 5022
rect 26012 5010 26292 5012
rect 26012 4958 26238 5010
rect 26290 4958 26292 5010
rect 26012 4956 26292 4958
rect 26012 4562 26068 4956
rect 26236 4946 26292 4956
rect 26012 4510 26014 4562
rect 26066 4510 26068 4562
rect 26012 4498 26068 4510
rect 26684 4562 26740 6636
rect 26684 4510 26686 4562
rect 26738 4510 26740 4562
rect 26684 4498 26740 4510
rect 25788 4340 25844 4350
rect 25788 4338 26404 4340
rect 25788 4286 25790 4338
rect 25842 4286 26404 4338
rect 25788 4284 26404 4286
rect 25788 4274 25844 4284
rect 26348 3778 26404 4284
rect 26348 3726 26350 3778
rect 26402 3726 26404 3778
rect 26348 3714 26404 3726
rect 26684 3780 26740 3790
rect 26796 3780 26852 7756
rect 26908 6468 26964 16716
rect 29708 16100 29764 16110
rect 28476 13748 28532 13758
rect 27804 8372 27860 8382
rect 27132 8148 27188 8158
rect 27132 8146 27524 8148
rect 27132 8094 27134 8146
rect 27186 8094 27524 8146
rect 27132 8092 27524 8094
rect 27132 8082 27188 8092
rect 27468 6914 27524 8092
rect 27804 8034 27860 8316
rect 27804 7982 27806 8034
rect 27858 7982 27860 8034
rect 27804 7812 27860 7982
rect 27804 7746 27860 7756
rect 27468 6862 27470 6914
rect 27522 6862 27524 6914
rect 27468 6850 27524 6862
rect 27804 6804 27860 6814
rect 27804 6710 27860 6748
rect 28140 6578 28196 6590
rect 28140 6526 28142 6578
rect 28194 6526 28196 6578
rect 26908 6466 27076 6468
rect 26908 6414 26910 6466
rect 26962 6414 27076 6466
rect 26908 6412 27076 6414
rect 26908 6402 26964 6412
rect 26908 6132 26964 6142
rect 26908 5122 26964 6076
rect 26908 5070 26910 5122
rect 26962 5070 26964 5122
rect 26908 5058 26964 5070
rect 27020 4338 27076 6412
rect 27804 5234 27860 5246
rect 27804 5182 27806 5234
rect 27858 5182 27860 5234
rect 27580 4452 27636 4462
rect 27580 4358 27636 4396
rect 27020 4286 27022 4338
rect 27074 4286 27076 4338
rect 27020 4274 27076 4286
rect 27468 4338 27524 4350
rect 27468 4286 27470 4338
rect 27522 4286 27524 4338
rect 26684 3778 26852 3780
rect 26684 3726 26686 3778
rect 26738 3726 26852 3778
rect 26684 3724 26852 3726
rect 27132 3780 27188 3790
rect 26684 3714 26740 3724
rect 26124 3444 26180 3454
rect 25676 3332 25732 3342
rect 25564 3330 25732 3332
rect 25564 3278 25678 3330
rect 25730 3278 25732 3330
rect 25564 3276 25732 3278
rect 25676 3266 25732 3276
rect 25340 3164 25620 3220
rect 24780 1026 24836 1036
rect 25564 800 25620 3164
rect 26124 800 26180 3388
rect 27132 3220 27188 3724
rect 27244 3556 27300 3566
rect 27244 3442 27300 3500
rect 27244 3390 27246 3442
rect 27298 3390 27300 3442
rect 27244 3378 27300 3390
rect 27468 3554 27524 4286
rect 27468 3502 27470 3554
rect 27522 3502 27524 3554
rect 27468 3444 27524 3502
rect 27468 3378 27524 3388
rect 27132 3164 27300 3220
rect 27244 800 27300 3164
rect 27804 800 27860 5182
rect 28140 3444 28196 6526
rect 28252 3556 28308 3566
rect 28252 3462 28308 3500
rect 28140 3378 28196 3388
rect 28476 3330 28532 13692
rect 28812 8034 28868 8046
rect 29596 8036 29652 8046
rect 28812 7982 28814 8034
rect 28866 7982 28868 8034
rect 28588 7362 28644 7374
rect 28588 7310 28590 7362
rect 28642 7310 28644 7362
rect 28588 6580 28644 7310
rect 28812 7364 28868 7982
rect 29260 8034 29652 8036
rect 29260 7982 29598 8034
rect 29650 7982 29652 8034
rect 29260 7980 29652 7982
rect 29148 7700 29204 7710
rect 29036 7364 29092 7374
rect 28812 7362 29092 7364
rect 28812 7310 29038 7362
rect 29090 7310 29092 7362
rect 28812 7308 29092 7310
rect 28588 6578 28756 6580
rect 28588 6526 28590 6578
rect 28642 6526 28756 6578
rect 28588 6524 28756 6526
rect 28588 6514 28644 6524
rect 28588 5794 28644 5806
rect 28588 5742 28590 5794
rect 28642 5742 28644 5794
rect 28588 4452 28644 5742
rect 28700 5122 28756 6524
rect 29036 6132 29092 7308
rect 29036 6066 29092 6076
rect 29148 6804 29204 7644
rect 29148 6130 29204 6748
rect 29148 6078 29150 6130
rect 29202 6078 29204 6130
rect 29148 6066 29204 6078
rect 28700 5070 28702 5122
rect 28754 5070 28756 5122
rect 28700 5058 28756 5070
rect 28924 5682 28980 5694
rect 28924 5630 28926 5682
rect 28978 5630 28980 5682
rect 28588 4386 28644 4396
rect 28588 4228 28644 4238
rect 28588 4134 28644 4172
rect 28476 3278 28478 3330
rect 28530 3278 28532 3330
rect 28476 3266 28532 3278
rect 28924 800 28980 5630
rect 29148 4338 29204 4350
rect 29148 4286 29150 4338
rect 29202 4286 29204 4338
rect 29148 4228 29204 4286
rect 29148 4162 29204 4172
rect 29260 3556 29316 7980
rect 29596 7970 29652 7980
rect 29596 7362 29652 7374
rect 29596 7310 29598 7362
rect 29650 7310 29652 7362
rect 29596 6580 29652 7310
rect 29484 6578 29652 6580
rect 29484 6526 29598 6578
rect 29650 6526 29652 6578
rect 29484 6524 29652 6526
rect 29484 5682 29540 6524
rect 29596 6514 29652 6524
rect 29484 5630 29486 5682
rect 29538 5630 29540 5682
rect 29484 5618 29540 5630
rect 29260 3490 29316 3500
rect 29484 3780 29540 3790
rect 29484 3554 29540 3724
rect 29484 3502 29486 3554
rect 29538 3502 29540 3554
rect 29484 3490 29540 3502
rect 29708 3330 29764 16044
rect 29932 12180 29988 12190
rect 29932 6578 29988 12124
rect 30716 9826 30772 9838
rect 30716 9774 30718 9826
rect 30770 9774 30772 9826
rect 30716 9604 30772 9774
rect 30716 8258 30772 9548
rect 30716 8206 30718 8258
rect 30770 8206 30772 8258
rect 30716 8194 30772 8206
rect 29932 6526 29934 6578
rect 29986 6526 29988 6578
rect 29932 6514 29988 6526
rect 30044 7362 30100 7374
rect 30044 7310 30046 7362
rect 30098 7310 30100 7362
rect 29932 5796 29988 5806
rect 29708 3278 29710 3330
rect 29762 3278 29764 3330
rect 29708 3266 29764 3278
rect 29820 5794 29988 5796
rect 29820 5742 29934 5794
rect 29986 5742 29988 5794
rect 29820 5740 29988 5742
rect 29820 980 29876 5740
rect 29932 5730 29988 5740
rect 29932 4898 29988 4910
rect 29932 4846 29934 4898
rect 29986 4846 29988 4898
rect 29932 4450 29988 4846
rect 29932 4398 29934 4450
rect 29986 4398 29988 4450
rect 29932 4386 29988 4398
rect 30044 3780 30100 7310
rect 30604 7364 30660 7374
rect 30940 7364 30996 7374
rect 31052 7364 31108 7374
rect 30604 7362 30884 7364
rect 30604 7310 30606 7362
rect 30658 7310 30884 7362
rect 30604 7308 30884 7310
rect 30604 7298 30660 7308
rect 30604 6692 30660 6702
rect 30492 6578 30548 6590
rect 30492 6526 30494 6578
rect 30546 6526 30548 6578
rect 30268 5010 30324 5022
rect 30268 4958 30270 5010
rect 30322 4958 30324 5010
rect 30268 3780 30324 4958
rect 30380 3780 30436 3790
rect 30268 3778 30436 3780
rect 30268 3726 30382 3778
rect 30434 3726 30436 3778
rect 30268 3724 30436 3726
rect 30044 3714 30100 3724
rect 30380 3714 30436 3724
rect 30492 3444 30548 6526
rect 30604 6132 30660 6636
rect 30604 5236 30660 6076
rect 30716 5236 30772 5246
rect 30604 5234 30772 5236
rect 30604 5182 30718 5234
rect 30770 5182 30772 5234
rect 30604 5180 30772 5182
rect 30716 5170 30772 5180
rect 30716 3780 30772 3790
rect 30828 3780 30884 7308
rect 30940 7362 31052 7364
rect 30940 7310 30942 7362
rect 30994 7310 31052 7362
rect 30940 7308 31052 7310
rect 30940 7298 30996 7308
rect 30940 6468 30996 6478
rect 30940 5906 30996 6412
rect 31052 6466 31108 7308
rect 31276 7140 31332 20132
rect 32956 17668 33012 17678
rect 31388 9716 31444 9726
rect 31388 9714 31892 9716
rect 31388 9662 31390 9714
rect 31442 9662 31892 9714
rect 31388 9660 31892 9662
rect 31388 9650 31444 9660
rect 31836 9266 31892 9660
rect 31836 9214 31838 9266
rect 31890 9214 31892 9266
rect 31836 9202 31892 9214
rect 32844 9604 32900 9614
rect 32844 9266 32900 9548
rect 32844 9214 32846 9266
rect 32898 9214 32900 9266
rect 32844 9202 32900 9214
rect 32172 9044 32228 9054
rect 32172 8950 32228 8988
rect 31500 8148 31556 8158
rect 31500 8146 32004 8148
rect 31500 8094 31502 8146
rect 31554 8094 32004 8146
rect 31500 8092 32004 8094
rect 31500 8082 31556 8092
rect 31948 7698 32004 8092
rect 31948 7646 31950 7698
rect 32002 7646 32004 7698
rect 31948 7634 32004 7646
rect 32284 7588 32340 7598
rect 32284 7494 32340 7532
rect 31276 7074 31332 7084
rect 31500 7362 31556 7374
rect 31500 7310 31502 7362
rect 31554 7310 31556 7362
rect 31052 6414 31054 6466
rect 31106 6414 31108 6466
rect 31052 6244 31108 6414
rect 31052 6178 31108 6188
rect 30940 5854 30942 5906
rect 30994 5854 30996 5906
rect 30940 5842 30996 5854
rect 31500 5908 31556 7310
rect 32844 7362 32900 7374
rect 32844 7310 32846 7362
rect 32898 7310 32900 7362
rect 32844 7252 32900 7310
rect 32844 7186 32900 7196
rect 32060 6802 32116 6814
rect 32060 6750 32062 6802
rect 32114 6750 32116 6802
rect 31612 6468 31668 6478
rect 32060 6468 32116 6750
rect 31612 6466 31780 6468
rect 31612 6414 31614 6466
rect 31666 6414 31780 6466
rect 31612 6412 31780 6414
rect 31612 6402 31668 6412
rect 31500 5842 31556 5852
rect 31612 5796 31668 5806
rect 31612 5702 31668 5740
rect 31500 5236 31556 5246
rect 30716 3778 30884 3780
rect 30716 3726 30718 3778
rect 30770 3726 30884 3778
rect 30716 3724 30884 3726
rect 30716 3714 30772 3724
rect 30492 3378 30548 3388
rect 30604 3556 30660 3566
rect 29484 924 29876 980
rect 29484 800 29540 924
rect 30604 800 30660 3500
rect 30828 1316 30884 3724
rect 31164 5234 31556 5236
rect 31164 5182 31502 5234
rect 31554 5182 31556 5234
rect 31164 5180 31556 5182
rect 30940 3444 30996 3454
rect 30940 3350 30996 3388
rect 30828 1250 30884 1260
rect 31164 800 31220 5180
rect 31500 5170 31556 5180
rect 31724 5012 31780 6412
rect 32060 6402 32116 6412
rect 32844 6132 32900 6142
rect 32956 6132 33012 17612
rect 33628 16772 33684 22428
rect 34860 22484 34916 116174
rect 35868 115892 35924 119200
rect 37436 117908 37492 119200
rect 37436 117852 37940 117908
rect 37884 116562 37940 117852
rect 37884 116510 37886 116562
rect 37938 116510 37940 116562
rect 37884 116498 37940 116510
rect 38892 116450 38948 116462
rect 38892 116398 38894 116450
rect 38946 116398 38948 116450
rect 38892 116340 38948 116398
rect 38892 116274 38948 116284
rect 39340 116340 39396 116350
rect 39340 116246 39396 116284
rect 40572 116004 40628 119200
rect 42140 117908 42196 119200
rect 42140 117852 42644 117908
rect 42588 116562 42644 117852
rect 45276 117572 45332 119200
rect 45276 117516 45780 117572
rect 42588 116510 42590 116562
rect 42642 116510 42644 116562
rect 42588 116498 42644 116510
rect 45724 116562 45780 117516
rect 45724 116510 45726 116562
rect 45778 116510 45780 116562
rect 45724 116498 45780 116510
rect 46844 116564 46900 119200
rect 49980 117236 50036 119200
rect 49980 117170 50036 117180
rect 50876 117236 50932 117246
rect 47068 116564 47124 116574
rect 46844 116562 47124 116564
rect 46844 116510 47070 116562
rect 47122 116510 47124 116562
rect 46844 116508 47124 116510
rect 47068 116498 47124 116508
rect 50876 116562 50932 117180
rect 50876 116510 50878 116562
rect 50930 116510 50932 116562
rect 50876 116498 50932 116510
rect 51548 116564 51604 119200
rect 54684 117012 54740 119200
rect 54684 116946 54740 116956
rect 55468 117012 55524 117022
rect 51548 116498 51604 116508
rect 53004 116564 53060 116574
rect 53004 116470 53060 116508
rect 55468 116562 55524 116956
rect 55468 116510 55470 116562
rect 55522 116510 55524 116562
rect 55468 116498 55524 116510
rect 56252 116564 56308 119200
rect 56252 116498 56308 116508
rect 57148 116564 57204 116574
rect 57148 116470 57204 116508
rect 43596 116452 43652 116462
rect 43596 116450 43764 116452
rect 43596 116398 43598 116450
rect 43650 116398 43764 116450
rect 43596 116396 43764 116398
rect 43596 116386 43652 116396
rect 43708 116228 43764 116396
rect 45276 116450 45332 116462
rect 45276 116398 45278 116450
rect 45330 116398 45332 116450
rect 44044 116228 44100 116238
rect 43708 116226 44100 116228
rect 43708 116174 44046 116226
rect 44098 116174 44100 116226
rect 43708 116172 44100 116174
rect 40572 115948 40740 116004
rect 35868 115826 35924 115836
rect 36764 115892 36820 115902
rect 35532 115778 35588 115790
rect 35532 115726 35534 115778
rect 35586 115726 35588 115778
rect 35196 115668 35252 115678
rect 35532 115668 35588 115726
rect 36092 115668 36148 115678
rect 35532 115666 36148 115668
rect 35532 115614 36094 115666
rect 36146 115614 36148 115666
rect 35532 115612 36148 115614
rect 35196 115574 35252 115612
rect 36092 115602 36148 115612
rect 36764 115554 36820 115836
rect 40684 115892 40740 115948
rect 40684 115826 40740 115836
rect 42252 115892 42308 115902
rect 40572 115778 40628 115790
rect 40572 115726 40574 115778
rect 40626 115726 40628 115778
rect 39676 115668 39732 115678
rect 39676 115574 39732 115612
rect 40236 115668 40292 115678
rect 40572 115668 40628 115726
rect 41580 115668 41636 115678
rect 40572 115666 41636 115668
rect 40572 115614 41582 115666
rect 41634 115614 41636 115666
rect 40572 115612 41636 115614
rect 40236 115574 40292 115612
rect 41580 115602 41636 115612
rect 36764 115502 36766 115554
rect 36818 115502 36820 115554
rect 36764 115490 36820 115502
rect 42252 115554 42308 115836
rect 42252 115502 42254 115554
rect 42306 115502 42308 115554
rect 42252 115490 42308 115502
rect 35196 115276 35460 115286
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35196 115210 35460 115220
rect 35196 113708 35460 113718
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35196 113642 35460 113652
rect 35196 112140 35460 112150
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35196 112074 35460 112084
rect 35196 110572 35460 110582
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35196 110506 35460 110516
rect 35196 109004 35460 109014
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35196 108938 35460 108948
rect 35196 107436 35460 107446
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35196 107370 35460 107380
rect 35196 105868 35460 105878
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35196 105802 35460 105812
rect 35196 104300 35460 104310
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35196 104234 35460 104244
rect 35196 102732 35460 102742
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35196 102666 35460 102676
rect 35196 101164 35460 101174
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35196 101098 35460 101108
rect 35196 99596 35460 99606
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35196 99530 35460 99540
rect 35196 98028 35460 98038
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35196 97962 35460 97972
rect 35196 96460 35460 96470
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35196 96394 35460 96404
rect 35196 94892 35460 94902
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35196 94826 35460 94836
rect 35196 93324 35460 93334
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35196 93258 35460 93268
rect 35196 91756 35460 91766
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35196 91690 35460 91700
rect 35196 90188 35460 90198
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35196 90122 35460 90132
rect 35196 88620 35460 88630
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35196 88554 35460 88564
rect 35196 87052 35460 87062
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35196 86986 35460 86996
rect 35196 85484 35460 85494
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35196 85418 35460 85428
rect 35196 83916 35460 83926
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35196 83850 35460 83860
rect 35196 82348 35460 82358
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35196 82282 35460 82292
rect 35196 80780 35460 80790
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35196 80714 35460 80724
rect 35196 79212 35460 79222
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35196 79146 35460 79156
rect 35196 77644 35460 77654
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35196 77578 35460 77588
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 43708 29428 43764 116172
rect 44044 116162 44100 116172
rect 45276 115890 45332 116398
rect 48076 116452 48132 116462
rect 48076 116358 48132 116396
rect 48748 116452 48804 116462
rect 50204 116452 50260 116462
rect 48748 116228 48804 116396
rect 49980 116450 50260 116452
rect 49980 116398 50206 116450
rect 50258 116398 50260 116450
rect 49980 116396 50260 116398
rect 48748 116226 48916 116228
rect 48748 116174 48750 116226
rect 48802 116174 48916 116226
rect 48748 116172 48916 116174
rect 48748 116162 48804 116172
rect 45276 115838 45278 115890
rect 45330 115838 45332 115890
rect 45276 115826 45332 115838
rect 44380 115668 44436 115678
rect 44380 115574 44436 115612
rect 45052 115668 45108 115678
rect 45052 115574 45108 115612
rect 48748 115668 48804 115678
rect 48748 115574 48804 115612
rect 48860 102508 48916 116172
rect 49980 115890 50036 116396
rect 50204 116386 50260 116396
rect 53788 116450 53844 116462
rect 53788 116398 53790 116450
rect 53842 116398 53844 116450
rect 50556 116060 50820 116070
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50556 115994 50820 116004
rect 49980 115838 49982 115890
rect 50034 115838 50036 115890
rect 49980 115826 50036 115838
rect 53788 115780 53844 116398
rect 54684 116450 54740 116462
rect 54684 116398 54686 116450
rect 54738 116398 54740 116450
rect 54684 115890 54740 116398
rect 57932 116450 57988 116462
rect 57932 116398 57934 116450
rect 57986 116398 57988 116450
rect 57932 116116 57988 116398
rect 57932 116050 57988 116060
rect 58380 116226 58436 116238
rect 58380 116174 58382 116226
rect 58434 116174 58436 116226
rect 58380 116116 58436 116174
rect 58380 116050 58436 116060
rect 54684 115838 54686 115890
rect 54738 115838 54740 115890
rect 54684 115826 54740 115838
rect 59388 115892 59444 119200
rect 60956 117908 61012 119200
rect 60956 117852 61460 117908
rect 61404 116562 61460 117852
rect 61404 116510 61406 116562
rect 61458 116510 61460 116562
rect 61404 116498 61460 116510
rect 62412 116452 62468 116462
rect 62412 116450 62916 116452
rect 62412 116398 62414 116450
rect 62466 116398 62916 116450
rect 62412 116396 62916 116398
rect 62412 116386 62468 116396
rect 62860 116226 62916 116396
rect 62860 116174 62862 116226
rect 62914 116174 62916 116226
rect 59388 115826 59444 115836
rect 60284 115892 60340 115902
rect 53676 115724 53788 115780
rect 49756 115668 49812 115678
rect 49756 115574 49812 115612
rect 50556 114492 50820 114502
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50556 114426 50820 114436
rect 50556 112924 50820 112934
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50556 112858 50820 112868
rect 50556 111356 50820 111366
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50556 111290 50820 111300
rect 50556 109788 50820 109798
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50556 109722 50820 109732
rect 50556 108220 50820 108230
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50556 108154 50820 108164
rect 50556 106652 50820 106662
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50556 106586 50820 106596
rect 50556 105084 50820 105094
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50556 105018 50820 105028
rect 50556 103516 50820 103526
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50556 103450 50820 103460
rect 53676 102508 53732 115724
rect 53788 115714 53844 115724
rect 55132 115780 55188 115790
rect 55132 115686 55188 115724
rect 59052 115778 59108 115790
rect 59052 115726 59054 115778
rect 59106 115726 59108 115778
rect 54460 115668 54516 115678
rect 54460 115574 54516 115612
rect 58716 115666 58772 115678
rect 58716 115614 58718 115666
rect 58770 115614 58772 115666
rect 53788 115556 53844 115566
rect 53788 115462 53844 115500
rect 58156 115556 58212 115566
rect 58156 115462 58212 115500
rect 58716 115556 58772 115614
rect 59052 115668 59108 115726
rect 59612 115668 59668 115678
rect 59052 115666 59668 115668
rect 59052 115614 59614 115666
rect 59666 115614 59668 115666
rect 59052 115612 59668 115614
rect 59612 115602 59668 115612
rect 58716 115490 58772 115500
rect 60284 115554 60340 115836
rect 60284 115502 60286 115554
rect 60338 115502 60340 115554
rect 60284 115490 60340 115502
rect 43708 29362 43764 29372
rect 48748 102452 48916 102508
rect 53564 102452 53732 102508
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 45276 27300 45332 27310
rect 41020 27076 41076 27086
rect 40012 26964 40068 26974
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 38556 23044 38612 23054
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34860 22418 34916 22428
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 33628 16706 33684 16716
rect 35084 19460 35140 19470
rect 35084 10052 35140 19404
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 37884 15428 37940 15438
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 36876 12404 36932 12414
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 36316 10052 36372 10062
rect 35084 9996 35476 10052
rect 33516 9938 33572 9950
rect 33516 9886 33518 9938
rect 33570 9886 33572 9938
rect 33516 9156 33572 9886
rect 33964 9604 34020 9614
rect 35196 9604 35252 9614
rect 33964 9510 34020 9548
rect 34860 9602 35252 9604
rect 34860 9550 35198 9602
rect 35250 9550 35252 9602
rect 34860 9548 35252 9550
rect 33516 9090 33572 9100
rect 34636 9156 34692 9166
rect 33740 9044 33796 9054
rect 33740 8950 33796 8988
rect 34076 9044 34132 9054
rect 34076 8950 34132 8988
rect 34524 9042 34580 9054
rect 34524 8990 34526 9042
rect 34578 8990 34580 9042
rect 33628 8370 33684 8382
rect 33628 8318 33630 8370
rect 33682 8318 33684 8370
rect 33628 8148 33684 8318
rect 34300 8148 34356 8158
rect 33628 8146 34356 8148
rect 33628 8094 34302 8146
rect 34354 8094 34356 8146
rect 33628 8092 34356 8094
rect 32844 6130 33012 6132
rect 32844 6078 32846 6130
rect 32898 6078 33012 6130
rect 32844 6076 33012 6078
rect 33068 7476 33124 7486
rect 32844 6066 32900 6076
rect 32620 5908 32676 5918
rect 32620 5814 32676 5852
rect 32060 5794 32116 5806
rect 32060 5742 32062 5794
rect 32114 5742 32116 5794
rect 32060 5684 32116 5742
rect 32060 5618 32116 5628
rect 33068 5572 33124 7420
rect 33516 7476 33572 7486
rect 33516 7382 33572 7420
rect 34188 7474 34244 7486
rect 34188 7422 34190 7474
rect 34242 7422 34244 7474
rect 34188 7252 34244 7422
rect 34188 7186 34244 7196
rect 34188 6580 34244 6590
rect 34188 6486 34244 6524
rect 34188 6020 34244 6030
rect 34188 5926 34244 5964
rect 33068 5234 33124 5516
rect 33068 5182 33070 5234
rect 33122 5182 33124 5234
rect 33068 5170 33124 5182
rect 33852 5906 33908 5918
rect 33852 5854 33854 5906
rect 33906 5854 33908 5906
rect 31724 4946 31780 4956
rect 32284 5122 32340 5134
rect 32284 5070 32286 5122
rect 32338 5070 32340 5122
rect 32060 4228 32116 4238
rect 32284 4228 32340 5070
rect 32060 4226 32340 4228
rect 32060 4174 32062 4226
rect 32114 4174 32340 4226
rect 32060 4172 32340 4174
rect 32508 4900 32564 4910
rect 31500 3444 31556 3454
rect 31500 3350 31556 3388
rect 32060 3444 32116 4172
rect 32060 3378 32116 3388
rect 32284 3780 32340 3790
rect 32284 800 32340 3724
rect 32508 3666 32564 4844
rect 33516 4900 33572 4910
rect 33516 4564 33572 4844
rect 33852 4900 33908 5854
rect 33852 4834 33908 4844
rect 33964 5908 34020 5918
rect 33516 4470 33572 4508
rect 32844 4340 32900 4350
rect 32844 4246 32900 4284
rect 32508 3614 32510 3666
rect 32562 3614 32564 3666
rect 32508 3602 32564 3614
rect 32844 3444 32900 3454
rect 32844 800 32900 3388
rect 33516 3444 33572 3454
rect 33516 3350 33572 3388
rect 33964 800 34020 5852
rect 34300 4338 34356 8092
rect 34524 7924 34580 8990
rect 34524 7858 34580 7868
rect 34636 7588 34692 9100
rect 34300 4286 34302 4338
rect 34354 4286 34356 4338
rect 34300 4274 34356 4286
rect 34412 7532 34692 7588
rect 34748 8146 34804 8158
rect 34748 8094 34750 8146
rect 34802 8094 34804 8146
rect 34748 7924 34804 8094
rect 34412 3554 34468 7532
rect 34636 7364 34692 7374
rect 34748 7364 34804 7868
rect 34636 7362 34804 7364
rect 34636 7310 34638 7362
rect 34690 7310 34804 7362
rect 34636 7308 34804 7310
rect 34636 7298 34692 7308
rect 34860 6692 34916 9548
rect 35196 9538 35252 9548
rect 35420 9266 35476 9996
rect 35420 9214 35422 9266
rect 35474 9214 35476 9266
rect 35420 9044 35476 9214
rect 35420 8978 35476 8988
rect 36204 9602 36260 9614
rect 36204 9550 36206 9602
rect 36258 9550 36260 9602
rect 35084 8932 35140 8942
rect 35084 8260 35140 8876
rect 35868 8932 35924 8942
rect 35868 8838 35924 8876
rect 35756 8818 35812 8830
rect 35756 8766 35758 8818
rect 35810 8766 35812 8818
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35084 8128 35140 8204
rect 35420 8034 35476 8046
rect 35420 7982 35422 8034
rect 35474 7982 35476 8034
rect 35420 7588 35476 7982
rect 35420 7522 35476 7532
rect 35308 7364 35364 7374
rect 35308 7270 35364 7308
rect 35756 7250 35812 8766
rect 36204 8428 36260 9550
rect 36316 8930 36372 9996
rect 36316 8878 36318 8930
rect 36370 8878 36372 8930
rect 36316 8818 36372 8878
rect 36316 8766 36318 8818
rect 36370 8766 36372 8818
rect 36316 8754 36372 8766
rect 36540 9716 36596 9726
rect 36204 8372 36372 8428
rect 36092 7476 36148 7514
rect 36092 7410 36148 7420
rect 35756 7198 35758 7250
rect 35810 7198 35812 7250
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35756 6804 35812 7198
rect 36092 7250 36148 7262
rect 36092 7198 36094 7250
rect 36146 7198 36148 7250
rect 34748 5908 34804 5918
rect 34748 5814 34804 5852
rect 34860 5124 34916 6636
rect 35532 6748 35812 6804
rect 35980 6804 36036 6814
rect 34972 6468 35028 6478
rect 34972 6130 35028 6412
rect 34972 6078 34974 6130
rect 35026 6078 35028 6130
rect 34972 6066 35028 6078
rect 35532 5908 35588 6748
rect 35980 6690 36036 6748
rect 35980 6638 35982 6690
rect 36034 6638 36036 6690
rect 35980 6626 36036 6638
rect 35532 5842 35588 5852
rect 35756 6578 35812 6590
rect 35756 6526 35758 6578
rect 35810 6526 35812 6578
rect 35084 5796 35140 5806
rect 35084 5702 35140 5740
rect 35644 5794 35700 5806
rect 35644 5742 35646 5794
rect 35698 5742 35700 5794
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35644 5236 35700 5742
rect 35756 5796 35812 6526
rect 35756 5730 35812 5740
rect 35644 5170 35700 5180
rect 34860 5058 34916 5068
rect 35980 5124 36036 5134
rect 35980 5030 36036 5068
rect 35196 5012 35252 5022
rect 35196 4918 35252 4956
rect 35644 4900 35700 4910
rect 34748 4228 34804 4238
rect 34412 3502 34414 3554
rect 34466 3502 34468 3554
rect 34412 3490 34468 3502
rect 34524 4226 34804 4228
rect 34524 4174 34750 4226
rect 34802 4174 34804 4226
rect 34524 4172 34804 4174
rect 34524 800 34580 4172
rect 34748 4162 34804 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35420 3444 35476 3454
rect 35420 3350 35476 3388
rect 35644 800 35700 4844
rect 36092 4900 36148 7198
rect 36204 6580 36260 6590
rect 36204 6486 36260 6524
rect 36092 4834 36148 4844
rect 36316 4788 36372 8372
rect 36428 8148 36484 8158
rect 36428 8054 36484 8092
rect 36540 6804 36596 9660
rect 36876 8036 36932 12348
rect 37772 10610 37828 10622
rect 37772 10558 37774 10610
rect 37826 10558 37828 10610
rect 36988 10276 37044 10286
rect 36988 9266 37044 10220
rect 36988 9214 36990 9266
rect 37042 9214 37044 9266
rect 36988 9202 37044 9214
rect 37660 9826 37716 9838
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 37660 9604 37716 9774
rect 37660 9044 37716 9548
rect 37660 8978 37716 8988
rect 37436 8930 37492 8942
rect 37436 8878 37438 8930
rect 37490 8878 37492 8930
rect 37436 8428 37492 8878
rect 37436 8372 37716 8428
rect 36876 7942 36932 7980
rect 37324 8148 37380 8158
rect 37324 7476 37380 8092
rect 37548 7476 37604 7486
rect 37324 7474 37604 7476
rect 37324 7422 37550 7474
rect 37602 7422 37604 7474
rect 37324 7420 37604 7422
rect 36540 6738 36596 6748
rect 36652 7362 36708 7374
rect 36652 7310 36654 7362
rect 36706 7310 36708 7362
rect 36428 6692 36484 6702
rect 36428 6598 36484 6636
rect 36652 6580 36708 7310
rect 36652 6514 36708 6524
rect 36988 7362 37044 7374
rect 36988 7310 36990 7362
rect 37042 7310 37044 7362
rect 36876 6468 36932 6478
rect 36876 6374 36932 6412
rect 36988 6132 37044 7310
rect 36988 6066 37044 6076
rect 35868 4226 35924 4238
rect 35868 4174 35870 4226
rect 35922 4174 35924 4226
rect 35868 4116 35924 4174
rect 35868 1428 35924 4060
rect 36316 3554 36372 4732
rect 36316 3502 36318 3554
rect 36370 3502 36372 3554
rect 36316 3490 36372 3502
rect 36764 6020 36820 6030
rect 35868 1362 35924 1372
rect 36204 3444 36260 3454
rect 36204 800 36260 3388
rect 36764 2436 36820 5964
rect 36876 5796 36932 5806
rect 36876 5234 36932 5740
rect 36876 5182 36878 5234
rect 36930 5182 36932 5234
rect 36876 5170 36932 5182
rect 36764 2370 36820 2380
rect 37324 800 37380 7420
rect 37548 7410 37604 7420
rect 37436 6692 37492 6702
rect 37436 6598 37492 6636
rect 37436 5460 37492 5470
rect 37436 3554 37492 5404
rect 37660 5236 37716 8372
rect 37772 8372 37828 10558
rect 37884 8820 37940 15372
rect 38556 10836 38612 22988
rect 38444 10780 38556 10836
rect 37996 10724 38052 10734
rect 37996 10722 38388 10724
rect 37996 10670 37998 10722
rect 38050 10670 38388 10722
rect 37996 10668 38388 10670
rect 37996 10658 38052 10668
rect 38108 10276 38164 10286
rect 37996 9044 38052 9054
rect 37996 8950 38052 8988
rect 37884 8764 38052 8820
rect 37884 8372 37940 8382
rect 37772 8370 37940 8372
rect 37772 8318 37886 8370
rect 37938 8318 37940 8370
rect 37772 8316 37940 8318
rect 37884 8306 37940 8316
rect 37772 8036 37828 8046
rect 37772 6690 37828 7980
rect 37884 7700 37940 7710
rect 37996 7700 38052 8764
rect 37884 7698 38052 7700
rect 37884 7646 37886 7698
rect 37938 7646 38052 7698
rect 37884 7644 38052 7646
rect 37884 7634 37940 7644
rect 38108 6804 38164 10220
rect 38332 9938 38388 10668
rect 38332 9886 38334 9938
rect 38386 9886 38388 9938
rect 38332 9874 38388 9886
rect 38220 8484 38276 8494
rect 38444 8484 38500 10780
rect 38556 10770 38612 10780
rect 39116 11170 39172 11182
rect 39116 11118 39118 11170
rect 39170 11118 39172 11170
rect 38780 10500 38836 10510
rect 39116 10500 39172 11118
rect 39564 11170 39620 11182
rect 39564 11118 39566 11170
rect 39618 11118 39620 11170
rect 39340 10836 39396 10846
rect 39340 10742 39396 10780
rect 38780 10498 39172 10500
rect 38780 10446 38782 10498
rect 38834 10446 39172 10498
rect 38780 10444 39172 10446
rect 38668 8932 38724 8942
rect 38668 8838 38724 8876
rect 38220 8482 38500 8484
rect 38220 8430 38222 8482
rect 38274 8430 38500 8482
rect 38220 8428 38500 8430
rect 38780 8428 38836 10444
rect 39228 8932 39284 8942
rect 38220 8418 38276 8428
rect 37772 6638 37774 6690
rect 37826 6638 37828 6690
rect 37772 6626 37828 6638
rect 37996 6748 38164 6804
rect 38668 8372 38836 8428
rect 39004 8596 39060 8606
rect 37772 6466 37828 6478
rect 37772 6414 37774 6466
rect 37826 6414 37828 6466
rect 37772 6018 37828 6414
rect 37996 6356 38052 6748
rect 38220 6692 38276 6702
rect 37772 5966 37774 6018
rect 37826 5966 37828 6018
rect 37772 5954 37828 5966
rect 37884 6300 38052 6356
rect 38108 6578 38164 6590
rect 38108 6526 38110 6578
rect 38162 6526 38164 6578
rect 37660 5170 37716 5180
rect 37884 5122 37940 6300
rect 38108 6132 38164 6526
rect 38108 6066 38164 6076
rect 37884 5070 37886 5122
rect 37938 5070 37940 5122
rect 37884 5058 37940 5070
rect 38220 5122 38276 6636
rect 38220 5070 38222 5122
rect 38274 5070 38276 5122
rect 37548 5010 37604 5022
rect 37548 4958 37550 5010
rect 37602 4958 37604 5010
rect 37548 4900 37604 4958
rect 37996 5012 38052 5022
rect 38220 5012 38276 5070
rect 37996 4918 38052 4956
rect 38108 4956 38220 5012
rect 37548 4834 37604 4844
rect 37996 4452 38052 4462
rect 38108 4452 38164 4956
rect 38220 4946 38276 4956
rect 38556 5908 38612 5918
rect 38668 5908 38724 8372
rect 38892 8258 38948 8270
rect 38892 8206 38894 8258
rect 38946 8206 38948 8258
rect 38892 8148 38948 8206
rect 38892 8082 38948 8092
rect 39004 8146 39060 8540
rect 39004 8094 39006 8146
rect 39058 8094 39060 8146
rect 39004 8082 39060 8094
rect 39228 7698 39284 8876
rect 39564 8428 39620 11118
rect 39900 10498 39956 10510
rect 39900 10446 39902 10498
rect 39954 10446 39956 10498
rect 39900 10052 39956 10446
rect 39900 9492 39956 9996
rect 39900 9426 39956 9436
rect 39228 7646 39230 7698
rect 39282 7646 39284 7698
rect 39228 7634 39284 7646
rect 39452 8372 39620 8428
rect 38780 7362 38836 7374
rect 38780 7310 38782 7362
rect 38834 7310 38836 7362
rect 38780 6692 38836 7310
rect 39004 7364 39060 7374
rect 38780 6626 38836 6636
rect 38892 6690 38948 6702
rect 38892 6638 38894 6690
rect 38946 6638 38948 6690
rect 38556 5906 38724 5908
rect 38556 5854 38558 5906
rect 38610 5854 38724 5906
rect 38556 5852 38724 5854
rect 38892 6580 38948 6638
rect 37996 4450 38164 4452
rect 37996 4398 37998 4450
rect 38050 4398 38164 4450
rect 37996 4396 38164 4398
rect 37996 4386 38052 4396
rect 38556 4340 38612 5852
rect 38668 5012 38724 5022
rect 38668 4918 38724 4956
rect 38892 4676 38948 6524
rect 39004 5010 39060 7308
rect 39004 4958 39006 5010
rect 39058 4958 39060 5010
rect 39004 4900 39060 4958
rect 39004 4834 39060 4844
rect 39116 6466 39172 6478
rect 39116 6414 39118 6466
rect 39170 6414 39172 6466
rect 38892 4620 39060 4676
rect 38668 4340 38724 4350
rect 38556 4338 38724 4340
rect 38556 4286 38670 4338
rect 38722 4286 38724 4338
rect 38556 4284 38724 4286
rect 38668 4228 38724 4284
rect 38668 4162 38724 4172
rect 37436 3502 37438 3554
rect 37490 3502 37492 3554
rect 37436 3490 37492 3502
rect 37884 3666 37940 3678
rect 37884 3614 37886 3666
rect 37938 3614 37940 3666
rect 37884 800 37940 3614
rect 39004 800 39060 4620
rect 39116 2996 39172 6414
rect 39452 6468 39508 8372
rect 39788 8036 39844 8046
rect 39564 8034 39844 8036
rect 39564 7982 39790 8034
rect 39842 7982 39844 8034
rect 39564 7980 39844 7982
rect 39564 7586 39620 7980
rect 39788 7970 39844 7980
rect 39564 7534 39566 7586
rect 39618 7534 39620 7586
rect 39564 7522 39620 7534
rect 39676 6580 39732 6590
rect 39676 6486 39732 6524
rect 40012 6578 40068 26908
rect 40236 25620 40292 25630
rect 40236 20188 40292 25564
rect 40124 20132 40292 20188
rect 40124 9268 40180 20132
rect 40908 10500 40964 10510
rect 40124 8370 40180 9212
rect 40460 9938 40516 9950
rect 40460 9886 40462 9938
rect 40514 9886 40516 9938
rect 40124 8318 40126 8370
rect 40178 8318 40180 8370
rect 40124 8306 40180 8318
rect 40236 8596 40292 8606
rect 40236 8428 40292 8540
rect 40460 8428 40516 9886
rect 40908 9938 40964 10444
rect 40908 9886 40910 9938
rect 40962 9886 40964 9938
rect 40908 9874 40964 9886
rect 40236 8372 40516 8428
rect 40796 8930 40852 8942
rect 40796 8878 40798 8930
rect 40850 8878 40852 8930
rect 40012 6526 40014 6578
rect 40066 6526 40068 6578
rect 40012 6514 40068 6526
rect 39452 6412 39620 6468
rect 39340 6132 39396 6142
rect 39340 6038 39396 6076
rect 39228 6018 39284 6030
rect 39228 5966 39230 6018
rect 39282 5966 39284 6018
rect 39228 5236 39284 5966
rect 39564 6020 39620 6412
rect 39452 5908 39508 5918
rect 39452 5814 39508 5852
rect 39564 5684 39620 5964
rect 39228 5170 39284 5180
rect 39340 5628 39620 5684
rect 40012 5794 40068 5806
rect 40012 5742 40014 5794
rect 40066 5742 40068 5794
rect 39340 4450 39396 5628
rect 40012 5348 40068 5742
rect 40012 5282 40068 5292
rect 39564 5010 39620 5022
rect 39564 4958 39566 5010
rect 39618 4958 39620 5010
rect 39340 4398 39342 4450
rect 39394 4398 39396 4450
rect 39452 4564 39508 4574
rect 39564 4564 39620 4958
rect 39508 4508 39620 4564
rect 39900 4898 39956 4910
rect 39900 4846 39902 4898
rect 39954 4846 39956 4898
rect 39452 4432 39508 4508
rect 39340 4386 39396 4398
rect 39676 4338 39732 4350
rect 39676 4286 39678 4338
rect 39730 4286 39732 4338
rect 39676 4004 39732 4286
rect 39900 4116 39956 4846
rect 40124 4900 40180 4910
rect 40124 4450 40180 4844
rect 40124 4398 40126 4450
rect 40178 4398 40180 4450
rect 40124 4386 40180 4398
rect 39900 4050 39956 4060
rect 39676 3938 39732 3948
rect 39116 2930 39172 2940
rect 39564 3666 39620 3678
rect 39564 3614 39566 3666
rect 39618 3614 39620 3666
rect 39564 800 39620 3614
rect 40236 3554 40292 8372
rect 40348 8148 40404 8158
rect 40348 8054 40404 8092
rect 40796 8146 40852 8878
rect 40796 8094 40798 8146
rect 40850 8094 40852 8146
rect 40460 7362 40516 7374
rect 40460 7310 40462 7362
rect 40514 7310 40516 7362
rect 40348 6580 40404 6590
rect 40348 5012 40404 6524
rect 40460 6244 40516 7310
rect 40572 6580 40628 6590
rect 40572 6486 40628 6524
rect 40796 6356 40852 8094
rect 40908 7362 40964 7374
rect 40908 7310 40910 7362
rect 40962 7310 40964 7362
rect 40908 6804 40964 7310
rect 40908 6738 40964 6748
rect 40908 6580 40964 6590
rect 41020 6580 41076 27020
rect 44716 22932 44772 22942
rect 43036 15876 43092 15886
rect 42700 10610 42756 10622
rect 42700 10558 42702 10610
rect 42754 10558 42756 10610
rect 41580 10500 41636 10510
rect 41468 9604 41524 9614
rect 40908 6578 41076 6580
rect 40908 6526 40910 6578
rect 40962 6526 41076 6578
rect 40908 6524 41076 6526
rect 41356 9602 41524 9604
rect 41356 9550 41470 9602
rect 41522 9550 41524 9602
rect 41356 9548 41524 9550
rect 41356 8596 41412 9548
rect 41468 9538 41524 9548
rect 41468 9268 41524 9278
rect 41580 9268 41636 10444
rect 42700 10500 42756 10558
rect 42700 10434 42756 10444
rect 42140 9602 42196 9614
rect 42588 9604 42644 9614
rect 42140 9550 42142 9602
rect 42194 9550 42196 9602
rect 41468 9266 41636 9268
rect 41468 9214 41470 9266
rect 41522 9214 41636 9266
rect 41468 9212 41636 9214
rect 41916 9268 41972 9278
rect 41468 9044 41524 9212
rect 41916 9174 41972 9212
rect 41468 8978 41524 8988
rect 41356 7364 41412 8540
rect 42140 8428 42196 9550
rect 42028 8372 42196 8428
rect 42476 9602 42644 9604
rect 42476 9550 42590 9602
rect 42642 9550 42644 9602
rect 42476 9548 42644 9550
rect 42476 8482 42532 9548
rect 42588 9538 42644 9548
rect 42588 9268 42644 9278
rect 43036 9268 43092 15820
rect 43260 11396 43316 11406
rect 43148 11172 43204 11182
rect 43148 9940 43204 11116
rect 43260 10052 43316 11340
rect 43372 10500 43428 10510
rect 43372 10498 43652 10500
rect 43372 10446 43374 10498
rect 43426 10446 43652 10498
rect 43372 10444 43652 10446
rect 43372 10434 43428 10444
rect 43260 9996 43428 10052
rect 43148 9938 43316 9940
rect 43148 9886 43150 9938
rect 43202 9886 43316 9938
rect 43148 9884 43316 9886
rect 43148 9874 43204 9884
rect 42588 9266 43092 9268
rect 42588 9214 42590 9266
rect 42642 9214 43038 9266
rect 43090 9214 43092 9266
rect 42588 9212 43092 9214
rect 42588 9202 42644 9212
rect 42476 8430 42478 8482
rect 42530 8430 42532 8482
rect 42476 8418 42532 8430
rect 41804 8036 41860 8046
rect 40908 6514 40964 6524
rect 41356 6468 41412 7308
rect 41468 8034 41860 8036
rect 41468 7982 41806 8034
rect 41858 7982 41860 8034
rect 41468 7980 41860 7982
rect 41468 6692 41524 7980
rect 41804 7970 41860 7980
rect 41580 7364 41636 7374
rect 41916 7364 41972 7374
rect 41580 7362 41748 7364
rect 41580 7310 41582 7362
rect 41634 7310 41748 7362
rect 41580 7308 41748 7310
rect 41580 7298 41636 7308
rect 41468 6636 41636 6692
rect 41468 6468 41524 6478
rect 41356 6466 41524 6468
rect 41356 6414 41470 6466
rect 41522 6414 41524 6466
rect 41356 6412 41524 6414
rect 41468 6402 41524 6412
rect 40796 6300 40964 6356
rect 40460 6178 40516 6188
rect 40460 6020 40516 6030
rect 40796 6020 40852 6030
rect 40460 5926 40516 5964
rect 40684 6018 40852 6020
rect 40684 5966 40798 6018
rect 40850 5966 40852 6018
rect 40684 5964 40852 5966
rect 40460 5236 40516 5246
rect 40460 5234 40628 5236
rect 40460 5182 40462 5234
rect 40514 5182 40628 5234
rect 40460 5180 40628 5182
rect 40460 5170 40516 5180
rect 40572 5012 40628 5180
rect 40348 4956 40516 5012
rect 40348 4340 40404 4350
rect 40348 4246 40404 4284
rect 40460 4228 40516 4956
rect 40572 4788 40628 4956
rect 40572 4722 40628 4732
rect 40572 4564 40628 4574
rect 40684 4564 40740 5964
rect 40796 5954 40852 5964
rect 40572 4562 40740 4564
rect 40572 4510 40574 4562
rect 40626 4510 40740 4562
rect 40572 4508 40740 4510
rect 40572 4498 40628 4508
rect 40684 4452 40740 4508
rect 40796 4564 40852 4602
rect 40796 4498 40852 4508
rect 40684 4386 40740 4396
rect 40796 4340 40852 4350
rect 40460 4172 40740 4228
rect 40236 3502 40238 3554
rect 40290 3502 40292 3554
rect 40236 3490 40292 3502
rect 40684 800 40740 4172
rect 40796 4116 40852 4284
rect 40796 4050 40852 4060
rect 40908 3556 40964 6300
rect 41356 6244 41412 6254
rect 41244 3668 41300 3678
rect 41132 3556 41188 3566
rect 40908 3554 41188 3556
rect 40908 3502 41134 3554
rect 41186 3502 41188 3554
rect 40908 3500 41188 3502
rect 41132 3490 41188 3500
rect 41244 800 41300 3612
rect 41356 3332 41412 6188
rect 41580 4788 41636 6636
rect 41692 6132 41748 7308
rect 41804 7362 41972 7364
rect 41804 7310 41918 7362
rect 41970 7310 41972 7362
rect 41804 7308 41972 7310
rect 41804 6692 41860 7308
rect 41916 7298 41972 7308
rect 41804 6578 41860 6636
rect 41804 6526 41806 6578
rect 41858 6526 41860 6578
rect 41804 6468 41860 6526
rect 41804 6402 41860 6412
rect 42028 6356 42084 8372
rect 42252 8036 42308 8046
rect 42252 7942 42308 7980
rect 42588 8034 42644 8046
rect 42588 7982 42590 8034
rect 42642 7982 42644 8034
rect 42588 7924 42644 7982
rect 42588 7858 42644 7868
rect 42812 7588 42868 7598
rect 42812 7494 42868 7532
rect 42476 7474 42532 7486
rect 42476 7422 42478 7474
rect 42530 7422 42532 7474
rect 42364 6690 42420 6702
rect 42364 6638 42366 6690
rect 42418 6638 42420 6690
rect 42028 6290 42084 6300
rect 42140 6580 42196 6590
rect 41916 6132 41972 6142
rect 41692 6130 41972 6132
rect 41692 6078 41918 6130
rect 41970 6078 41972 6130
rect 41692 6076 41972 6078
rect 41916 5796 41972 6076
rect 41916 5730 41972 5740
rect 41580 4722 41636 4732
rect 41692 4228 41748 4238
rect 41692 4134 41748 4172
rect 42140 4116 42196 6524
rect 42364 5908 42420 6638
rect 42476 6692 42532 7422
rect 42476 6626 42532 6636
rect 42924 6690 42980 9212
rect 43036 9202 43092 9212
rect 43036 8596 43092 8606
rect 43036 8370 43092 8540
rect 43036 8318 43038 8370
rect 43090 8318 43092 8370
rect 43036 8306 43092 8318
rect 43148 8482 43204 8494
rect 43148 8430 43150 8482
rect 43202 8430 43204 8482
rect 42924 6638 42926 6690
rect 42978 6638 42980 6690
rect 42588 6578 42644 6590
rect 42588 6526 42590 6578
rect 42642 6526 42644 6578
rect 42252 5906 42420 5908
rect 42252 5854 42366 5906
rect 42418 5854 42420 5906
rect 42252 5852 42420 5854
rect 42252 4340 42308 5852
rect 42364 5842 42420 5852
rect 42476 6020 42532 6030
rect 42588 6020 42644 6526
rect 42812 6578 42868 6590
rect 42812 6526 42814 6578
rect 42866 6526 42868 6578
rect 42476 6018 42644 6020
rect 42476 5966 42478 6018
rect 42530 5966 42644 6018
rect 42476 5964 42644 5966
rect 42700 6356 42756 6366
rect 42700 6018 42756 6300
rect 42812 6244 42868 6526
rect 42812 6178 42868 6188
rect 42700 5966 42702 6018
rect 42754 5966 42756 6018
rect 42364 4452 42420 4462
rect 42476 4452 42532 5964
rect 42700 5954 42756 5966
rect 42924 5908 42980 6638
rect 42812 5906 42980 5908
rect 42812 5854 42926 5906
rect 42978 5854 42980 5906
rect 42812 5852 42980 5854
rect 42812 5684 42868 5852
rect 42924 5842 42980 5852
rect 43036 7924 43092 7934
rect 42588 5236 42644 5246
rect 42588 5142 42644 5180
rect 42420 4396 42532 4452
rect 42364 4358 42420 4396
rect 42252 4208 42308 4284
rect 42588 4340 42644 4350
rect 42140 4060 42420 4116
rect 41804 3668 41860 3678
rect 41804 3574 41860 3612
rect 41356 3266 41412 3276
rect 42364 800 42420 4060
rect 42588 3780 42644 4284
rect 42812 4338 42868 5628
rect 43036 5012 43092 7868
rect 43036 4946 43092 4956
rect 42812 4286 42814 4338
rect 42866 4286 42868 4338
rect 42812 4274 42868 4286
rect 43148 4340 43204 8430
rect 43260 7476 43316 9884
rect 43372 8428 43428 9996
rect 43596 9940 43652 10444
rect 43596 9884 43708 9940
rect 43652 9726 43708 9884
rect 43652 9714 43764 9726
rect 43652 9662 43710 9714
rect 43762 9662 43764 9714
rect 43652 9660 43764 9662
rect 43708 9650 43764 9660
rect 44044 9716 44100 9726
rect 44044 9714 44660 9716
rect 44044 9662 44046 9714
rect 44098 9662 44660 9714
rect 44044 9660 44660 9662
rect 44044 9650 44100 9660
rect 43484 9492 43540 9502
rect 43484 9266 43540 9436
rect 43484 9214 43486 9266
rect 43538 9214 43540 9266
rect 43484 9044 43540 9214
rect 44604 9266 44660 9660
rect 44604 9214 44606 9266
rect 44658 9214 44660 9266
rect 44604 9202 44660 9214
rect 43484 8978 43540 8988
rect 43932 9044 43988 9054
rect 43372 8372 43540 8428
rect 43372 7476 43428 7486
rect 43260 7474 43428 7476
rect 43260 7422 43374 7474
rect 43426 7422 43428 7474
rect 43260 7420 43428 7422
rect 43260 5124 43316 7420
rect 43372 7410 43428 7420
rect 43372 6692 43428 6702
rect 43484 6692 43540 8372
rect 43932 8370 43988 8988
rect 44380 9044 44436 9054
rect 43932 8318 43934 8370
rect 43986 8318 43988 8370
rect 43932 8306 43988 8318
rect 44044 8930 44100 8942
rect 44044 8878 44046 8930
rect 44098 8878 44100 8930
rect 44044 8260 44100 8878
rect 44044 8194 44100 8204
rect 43708 8034 43764 8046
rect 43708 7982 43710 8034
rect 43762 7982 43764 8034
rect 43708 7812 43764 7982
rect 43820 8036 43876 8046
rect 43820 8034 44324 8036
rect 43820 7982 43822 8034
rect 43874 7982 44324 8034
rect 43820 7980 44324 7982
rect 43820 7970 43876 7980
rect 43708 7746 43764 7756
rect 43932 7812 43988 7822
rect 43372 6690 43540 6692
rect 43372 6638 43374 6690
rect 43426 6638 43540 6690
rect 43372 6636 43540 6638
rect 43372 6626 43428 6636
rect 43820 6468 43876 6478
rect 43820 6374 43876 6412
rect 43932 6244 43988 7756
rect 44156 7588 44212 7598
rect 44156 7494 44212 7532
rect 43820 6188 43988 6244
rect 44044 6580 44100 6590
rect 43260 4992 43316 5068
rect 43372 5682 43428 5694
rect 43372 5630 43374 5682
rect 43426 5630 43428 5682
rect 43372 4900 43428 5630
rect 43372 4834 43428 4844
rect 43260 4452 43316 4462
rect 43260 4358 43316 4396
rect 43148 4274 43204 4284
rect 42588 3714 42644 3724
rect 43148 3666 43204 3678
rect 43148 3614 43150 3666
rect 43202 3614 43204 3666
rect 43148 980 43204 3614
rect 43820 3332 43876 6188
rect 43932 5122 43988 5134
rect 43932 5070 43934 5122
rect 43986 5070 43988 5122
rect 43932 5012 43988 5070
rect 43932 4946 43988 4956
rect 44044 3554 44100 6524
rect 44268 6244 44324 7980
rect 44380 6578 44436 8988
rect 44380 6526 44382 6578
rect 44434 6526 44436 6578
rect 44380 6514 44436 6526
rect 44604 6690 44660 6702
rect 44604 6638 44606 6690
rect 44658 6638 44660 6690
rect 44604 6468 44660 6638
rect 44604 6402 44660 6412
rect 44268 6188 44660 6244
rect 44156 6020 44212 6030
rect 44156 5926 44212 5964
rect 44604 6018 44660 6188
rect 44604 5966 44606 6018
rect 44658 5966 44660 6018
rect 44604 5954 44660 5966
rect 44380 5010 44436 5022
rect 44380 4958 44382 5010
rect 44434 4958 44436 5010
rect 44380 4788 44436 4958
rect 44716 5010 44772 22876
rect 44940 10836 44996 10846
rect 44828 9602 44884 9614
rect 44828 9550 44830 9602
rect 44882 9550 44884 9602
rect 44828 8596 44884 9550
rect 44940 9042 44996 10780
rect 45276 10836 45332 27244
rect 45276 10770 45332 10780
rect 45724 27188 45780 27198
rect 44940 8990 44942 9042
rect 44994 8990 44996 9042
rect 44940 8978 44996 8990
rect 45052 10724 45108 10734
rect 44828 8530 44884 8540
rect 44828 8034 44884 8046
rect 44828 7982 44830 8034
rect 44882 7982 44884 8034
rect 44828 7812 44884 7982
rect 44828 7746 44884 7756
rect 45052 8036 45108 10668
rect 45724 10612 45780 27132
rect 48636 23828 48692 23838
rect 46956 23716 47012 23726
rect 46284 21364 46340 21374
rect 45724 10546 45780 10556
rect 46172 11620 46228 11630
rect 45500 10500 45556 10510
rect 45388 10498 45556 10500
rect 45388 10446 45502 10498
rect 45554 10446 45556 10498
rect 45388 10444 45556 10446
rect 45388 9156 45444 10444
rect 45500 10434 45556 10444
rect 46060 10500 46116 10510
rect 46060 10406 46116 10444
rect 45612 9826 45668 9838
rect 45612 9774 45614 9826
rect 45666 9774 45668 9826
rect 45500 9156 45556 9166
rect 45388 9154 45556 9156
rect 45388 9102 45502 9154
rect 45554 9102 45556 9154
rect 45388 9100 45556 9102
rect 45388 8428 45444 9100
rect 45500 9090 45556 9100
rect 45052 7476 45108 7980
rect 44828 7420 45108 7476
rect 45164 8372 45444 8428
rect 45500 8596 45556 8606
rect 45612 8596 45668 9774
rect 45836 9602 45892 9614
rect 46172 9604 46228 11564
rect 45836 9550 45838 9602
rect 45890 9550 45892 9602
rect 45724 9380 45780 9390
rect 45724 9042 45780 9324
rect 45836 9268 45892 9550
rect 45836 9202 45892 9212
rect 46060 9548 46228 9604
rect 45724 8990 45726 9042
rect 45778 8990 45780 9042
rect 45724 8978 45780 8990
rect 45556 8540 45668 8596
rect 45724 8820 45780 8830
rect 44828 6018 44884 7420
rect 45164 6356 45220 8372
rect 45500 8258 45556 8540
rect 45724 8428 45780 8764
rect 46060 8428 46116 9548
rect 45500 8206 45502 8258
rect 45554 8206 45556 8258
rect 45500 8194 45556 8206
rect 45612 8372 45780 8428
rect 45948 8372 46116 8428
rect 46172 9380 46228 9390
rect 45612 6916 45668 8372
rect 44828 5966 44830 6018
rect 44882 5966 44884 6018
rect 44828 5954 44884 5966
rect 44940 6300 45220 6356
rect 45500 6860 45668 6916
rect 45724 8260 45780 8270
rect 45724 8036 45780 8204
rect 44716 4958 44718 5010
rect 44770 4958 44772 5010
rect 44716 4946 44772 4958
rect 44044 3502 44046 3554
rect 44098 3502 44100 3554
rect 44044 3490 44100 3502
rect 44268 4226 44324 4238
rect 44268 4174 44270 4226
rect 44322 4174 44324 4226
rect 43820 3276 44100 3332
rect 42924 924 43204 980
rect 42924 800 42980 924
rect 44044 800 44100 3276
rect 44268 2212 44324 4174
rect 44380 4228 44436 4732
rect 44940 4338 44996 6300
rect 45276 5906 45332 5918
rect 45276 5854 45278 5906
rect 45330 5854 45332 5906
rect 45052 5794 45108 5806
rect 45052 5742 45054 5794
rect 45106 5742 45108 5794
rect 45052 5236 45108 5742
rect 45276 5796 45332 5854
rect 45276 5730 45332 5740
rect 45500 5796 45556 6860
rect 45612 6692 45668 6702
rect 45612 6598 45668 6636
rect 45500 5730 45556 5740
rect 45052 5170 45108 5180
rect 44940 4286 44942 4338
rect 44994 4286 44996 4338
rect 44940 4274 44996 4286
rect 45388 5122 45444 5134
rect 45388 5070 45390 5122
rect 45442 5070 45444 5122
rect 45388 4340 45444 5070
rect 45388 4274 45444 4284
rect 44380 4162 44436 4172
rect 45500 4226 45556 4238
rect 45500 4174 45502 4226
rect 45554 4174 45556 4226
rect 45500 3556 45556 4174
rect 45500 3490 45556 3500
rect 45388 3444 45444 3454
rect 45388 3350 45444 3388
rect 44268 2156 44660 2212
rect 44604 800 44660 2156
rect 45724 800 45780 7980
rect 45836 8034 45892 8046
rect 45836 7982 45838 8034
rect 45890 7982 45892 8034
rect 45836 7140 45892 7982
rect 45836 7074 45892 7084
rect 45948 6914 46004 8372
rect 46172 7364 46228 9324
rect 46284 7588 46340 21308
rect 46844 17556 46900 17566
rect 46620 11172 46676 11182
rect 46396 10836 46452 10846
rect 46396 10742 46452 10780
rect 46620 10836 46676 11116
rect 46620 10770 46676 10780
rect 46620 10612 46676 10622
rect 46508 9156 46564 9166
rect 46508 9062 46564 9100
rect 46396 8146 46452 8158
rect 46396 8094 46398 8146
rect 46450 8094 46452 8146
rect 46396 8036 46452 8094
rect 46396 7970 46452 7980
rect 46284 7532 46452 7588
rect 46172 7298 46228 7308
rect 46284 7362 46340 7374
rect 46284 7310 46286 7362
rect 46338 7310 46340 7362
rect 45948 6862 45950 6914
rect 46002 6862 46004 6914
rect 45948 6850 46004 6862
rect 46172 6692 46228 6702
rect 46060 6356 46116 6366
rect 45948 6244 46004 6254
rect 45948 5348 46004 6188
rect 46060 6130 46116 6300
rect 46060 6078 46062 6130
rect 46114 6078 46116 6130
rect 46060 6066 46116 6078
rect 46172 6020 46228 6636
rect 46284 6580 46340 7310
rect 46396 6692 46452 7532
rect 46396 6626 46452 6636
rect 46284 6514 46340 6524
rect 46508 6580 46564 6590
rect 46508 6486 46564 6524
rect 46172 5954 46228 5964
rect 46396 6468 46452 6478
rect 45948 5216 46004 5292
rect 46284 5908 46340 5918
rect 46284 5346 46340 5852
rect 46284 5294 46286 5346
rect 46338 5294 46340 5346
rect 46284 5282 46340 5294
rect 46172 4898 46228 4910
rect 46172 4846 46174 4898
rect 46226 4846 46228 4898
rect 46172 3780 46228 4846
rect 46172 3714 46228 3724
rect 46060 3556 46116 3566
rect 46396 3556 46452 6412
rect 46620 6132 46676 10556
rect 46732 10500 46788 10510
rect 46732 9826 46788 10444
rect 46732 9774 46734 9826
rect 46786 9774 46788 9826
rect 46732 9762 46788 9774
rect 46844 9604 46900 17500
rect 46956 11620 47012 23660
rect 47964 17108 48020 17118
rect 47012 11564 47236 11620
rect 46956 11488 47012 11564
rect 47180 11506 47236 11564
rect 47180 11454 47182 11506
rect 47234 11454 47236 11506
rect 47180 11442 47236 11454
rect 47628 11172 47684 11182
rect 47292 11170 47684 11172
rect 47292 11118 47630 11170
rect 47682 11118 47684 11170
rect 47292 11116 47684 11118
rect 47292 10724 47348 11116
rect 47628 11106 47684 11116
rect 47628 10724 47684 10734
rect 46732 9548 46900 9604
rect 47068 10668 47348 10724
rect 47404 10722 47684 10724
rect 47404 10670 47630 10722
rect 47682 10670 47684 10722
rect 47404 10668 47684 10670
rect 46732 8146 46788 9548
rect 46844 9268 46900 9278
rect 46844 9174 46900 9212
rect 47068 8428 47124 10668
rect 46732 8094 46734 8146
rect 46786 8094 46788 8146
rect 46732 8082 46788 8094
rect 46956 8372 47124 8428
rect 47180 10498 47236 10510
rect 47180 10446 47182 10498
rect 47234 10446 47236 10498
rect 47180 9156 47236 10446
rect 47404 9938 47460 10668
rect 47628 10658 47684 10668
rect 47852 10612 47908 10622
rect 47404 9886 47406 9938
rect 47458 9886 47460 9938
rect 47404 9874 47460 9886
rect 47740 10610 47908 10612
rect 47740 10558 47854 10610
rect 47906 10558 47908 10610
rect 47740 10556 47908 10558
rect 47516 9268 47572 9278
rect 47740 9268 47796 10556
rect 47852 10546 47908 10556
rect 47516 9266 47796 9268
rect 47516 9214 47518 9266
rect 47570 9214 47796 9266
rect 47516 9212 47796 9214
rect 47852 10388 47908 10398
rect 47516 9202 47572 9212
rect 46956 7476 47012 8372
rect 46956 7382 47012 7420
rect 46732 7364 46788 7374
rect 46732 6690 46788 7308
rect 46732 6638 46734 6690
rect 46786 6638 46788 6690
rect 46732 6626 46788 6638
rect 46844 6132 46900 6142
rect 46620 6130 46900 6132
rect 46620 6078 46846 6130
rect 46898 6078 46900 6130
rect 46620 6076 46900 6078
rect 46844 6066 46900 6076
rect 46620 5906 46676 5918
rect 46620 5854 46622 5906
rect 46674 5854 46676 5906
rect 46620 5684 46676 5854
rect 46620 5618 46676 5628
rect 47180 4228 47236 9100
rect 47852 9042 47908 10332
rect 47852 8990 47854 9042
rect 47906 8990 47908 9042
rect 47852 8978 47908 8990
rect 47964 8428 48020 17052
rect 47404 8372 48020 8428
rect 48076 11170 48132 11182
rect 48076 11118 48078 11170
rect 48130 11118 48132 11170
rect 47292 8146 47348 8158
rect 47292 8094 47294 8146
rect 47346 8094 47348 8146
rect 47292 7924 47348 8094
rect 47292 7858 47348 7868
rect 47292 7700 47348 7710
rect 47404 7700 47460 8372
rect 47292 7698 47460 7700
rect 47292 7646 47294 7698
rect 47346 7646 47460 7698
rect 47292 7644 47460 7646
rect 47628 8034 47684 8046
rect 47628 7982 47630 8034
rect 47682 7982 47684 8034
rect 47292 7634 47348 7644
rect 47628 6804 47684 7982
rect 47852 7474 47908 7486
rect 47852 7422 47854 7474
rect 47906 7422 47908 7474
rect 47852 7252 47908 7422
rect 47852 7186 47908 7196
rect 48076 6804 48132 11118
rect 48636 10836 48692 23772
rect 48748 21028 48804 102452
rect 50556 101948 50820 101958
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50556 101882 50820 101892
rect 50556 100380 50820 100390
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50556 100314 50820 100324
rect 50556 98812 50820 98822
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50556 98746 50820 98756
rect 50556 97244 50820 97254
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50556 97178 50820 97188
rect 50556 95676 50820 95686
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50556 95610 50820 95620
rect 50556 94108 50820 94118
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50556 94042 50820 94052
rect 50556 92540 50820 92550
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50556 92474 50820 92484
rect 50556 90972 50820 90982
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50556 90906 50820 90916
rect 50556 89404 50820 89414
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50556 89338 50820 89348
rect 50556 87836 50820 87846
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50556 87770 50820 87780
rect 50556 86268 50820 86278
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50556 86202 50820 86212
rect 50556 84700 50820 84710
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50556 84634 50820 84644
rect 50556 83132 50820 83142
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50556 83066 50820 83076
rect 50556 81564 50820 81574
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50556 81498 50820 81508
rect 50556 79996 50820 80006
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50556 79930 50820 79940
rect 50556 78428 50820 78438
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50556 78362 50820 78372
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 48748 20962 48804 20972
rect 49196 30324 49252 30334
rect 49196 20188 49252 30268
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 52780 25508 52836 25518
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 49196 20132 49364 20188
rect 48972 16996 49028 17006
rect 48748 11172 48804 11182
rect 48748 11170 48916 11172
rect 48748 11118 48750 11170
rect 48802 11118 48916 11170
rect 48748 11116 48916 11118
rect 48748 11106 48804 11116
rect 48748 10836 48804 10846
rect 48636 10834 48804 10836
rect 48636 10782 48750 10834
rect 48802 10782 48804 10834
rect 48636 10780 48804 10782
rect 48636 10388 48692 10780
rect 48748 10770 48804 10780
rect 48636 10322 48692 10332
rect 48300 9156 48356 9166
rect 47628 6738 47684 6748
rect 47852 6748 48132 6804
rect 48188 8370 48244 8382
rect 48188 8318 48190 8370
rect 48242 8318 48244 8370
rect 47740 6692 47796 6702
rect 47740 6580 47796 6636
rect 47628 6578 47796 6580
rect 47628 6526 47742 6578
rect 47794 6526 47796 6578
rect 47628 6524 47796 6526
rect 47628 6244 47684 6524
rect 47740 6514 47796 6524
rect 47628 6178 47684 6188
rect 47740 6130 47796 6142
rect 47740 6078 47742 6130
rect 47794 6078 47796 6130
rect 47628 6020 47684 6030
rect 47628 5926 47684 5964
rect 47404 5908 47460 5918
rect 47404 5814 47460 5852
rect 47404 5236 47460 5246
rect 47404 5234 47572 5236
rect 47404 5182 47406 5234
rect 47458 5182 47572 5234
rect 47404 5180 47572 5182
rect 47404 5170 47460 5180
rect 47180 4172 47460 4228
rect 46060 3554 46452 3556
rect 46060 3502 46062 3554
rect 46114 3502 46452 3554
rect 46060 3500 46452 3502
rect 46844 3556 46900 3566
rect 46060 3490 46116 3500
rect 46844 3462 46900 3500
rect 46284 3332 46340 3342
rect 46284 800 46340 3276
rect 47404 800 47460 4172
rect 47516 1764 47572 5180
rect 47628 4452 47684 4462
rect 47740 4452 47796 6078
rect 47852 5684 47908 6748
rect 48076 6578 48132 6590
rect 48076 6526 48078 6578
rect 48130 6526 48132 6578
rect 48076 6132 48132 6526
rect 48188 6468 48244 8318
rect 48188 6402 48244 6412
rect 48076 6066 48132 6076
rect 47964 5906 48020 5918
rect 47964 5854 47966 5906
rect 48018 5854 48020 5906
rect 47964 5796 48020 5854
rect 47964 5730 48020 5740
rect 47852 5618 47908 5628
rect 48300 5460 48356 9100
rect 48636 9156 48692 9166
rect 48636 9062 48692 9100
rect 48412 9042 48468 9054
rect 48412 8990 48414 9042
rect 48466 8990 48468 9042
rect 48412 7364 48468 8990
rect 48860 8428 48916 11116
rect 48972 9268 49028 16940
rect 48972 9202 49028 9212
rect 49084 10052 49140 10062
rect 48412 7270 48468 7308
rect 48636 8372 48916 8428
rect 48636 7252 48692 8372
rect 48636 6578 48692 7196
rect 48636 6526 48638 6578
rect 48690 6526 48692 6578
rect 48636 6514 48692 6526
rect 48748 7476 48804 7486
rect 48076 5404 48356 5460
rect 48076 5122 48132 5404
rect 48076 5070 48078 5122
rect 48130 5070 48132 5122
rect 48076 5058 48132 5070
rect 47628 4450 47796 4452
rect 47628 4398 47630 4450
rect 47682 4398 47796 4450
rect 47628 4396 47796 4398
rect 47628 4386 47684 4396
rect 48412 4340 48468 4350
rect 48412 4246 48468 4284
rect 47740 3444 47796 3454
rect 48748 3444 48804 7420
rect 48972 6580 49028 6590
rect 48972 6356 49028 6524
rect 48972 6290 49028 6300
rect 48860 6020 48916 6030
rect 48860 5926 48916 5964
rect 49084 5460 49140 9996
rect 48860 5012 48916 5022
rect 48860 4918 48916 4956
rect 49084 3666 49140 5404
rect 49196 5012 49252 5022
rect 49308 5012 49364 20132
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 51548 12516 51604 12526
rect 51100 11284 51156 11294
rect 51100 11190 51156 11228
rect 51324 11284 51380 11294
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 51100 10836 51156 10846
rect 50876 10612 50932 10622
rect 49868 10500 49924 10510
rect 49868 10406 49924 10444
rect 50652 10500 50708 10510
rect 50876 10500 50932 10556
rect 50652 10498 50932 10500
rect 50652 10446 50654 10498
rect 50706 10446 50932 10498
rect 50652 10444 50932 10446
rect 50652 10434 50708 10444
rect 49532 9938 49588 9950
rect 49532 9886 49534 9938
rect 49586 9886 49588 9938
rect 49532 9156 49588 9886
rect 50876 9938 50932 10444
rect 50876 9886 50878 9938
rect 50930 9886 50932 9938
rect 50428 9714 50484 9726
rect 50428 9662 50430 9714
rect 50482 9662 50484 9714
rect 49532 9090 49588 9100
rect 50092 9602 50148 9614
rect 50092 9550 50094 9602
rect 50146 9550 50148 9602
rect 49980 9044 50036 9054
rect 49756 7364 49812 7374
rect 49756 6690 49812 7308
rect 49756 6638 49758 6690
rect 49810 6638 49812 6690
rect 49756 6626 49812 6638
rect 49644 6578 49700 6590
rect 49644 6526 49646 6578
rect 49698 6526 49700 6578
rect 49644 6468 49700 6526
rect 49644 6402 49700 6412
rect 49980 6020 50036 8988
rect 50092 8428 50148 9550
rect 50316 9044 50372 9054
rect 50316 8950 50372 8988
rect 50092 8372 50372 8428
rect 50316 8370 50372 8372
rect 50316 8318 50318 8370
rect 50370 8318 50372 8370
rect 50316 8306 50372 8318
rect 50428 7588 50484 9662
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50428 7532 50820 7588
rect 50428 7028 50484 7038
rect 50428 6914 50484 6972
rect 50428 6862 50430 6914
rect 50482 6862 50484 6914
rect 50428 6850 50484 6862
rect 50764 6690 50820 7532
rect 50764 6638 50766 6690
rect 50818 6638 50820 6690
rect 50764 6626 50820 6638
rect 50876 6692 50932 9886
rect 50988 8258 51044 8270
rect 50988 8206 50990 8258
rect 51042 8206 51044 8258
rect 50988 7924 51044 8206
rect 50988 7858 51044 7868
rect 51100 7586 51156 10780
rect 51212 10498 51268 10510
rect 51212 10446 51214 10498
rect 51266 10446 51268 10498
rect 51212 10052 51268 10446
rect 51212 9986 51268 9996
rect 51324 8428 51380 11228
rect 51548 10388 51604 12460
rect 52780 12404 52836 25452
rect 52108 12402 52836 12404
rect 52108 12350 52782 12402
rect 52834 12350 52836 12402
rect 52108 12348 52836 12350
rect 51996 11844 52052 11854
rect 51996 11508 52052 11788
rect 51772 11506 52052 11508
rect 51772 11454 51998 11506
rect 52050 11454 52052 11506
rect 51772 11452 52052 11454
rect 51660 11172 51716 11182
rect 51660 11078 51716 11116
rect 51772 10722 51828 11452
rect 51996 11442 52052 11452
rect 51772 10670 51774 10722
rect 51826 10670 51828 10722
rect 51772 10658 51828 10670
rect 51884 10612 51940 10622
rect 51660 10388 51716 10398
rect 51548 10386 51716 10388
rect 51548 10334 51662 10386
rect 51714 10334 51716 10386
rect 51548 10332 51716 10334
rect 51100 7534 51102 7586
rect 51154 7534 51156 7586
rect 51100 7522 51156 7534
rect 51212 8372 51380 8428
rect 51436 9826 51492 9838
rect 51436 9774 51438 9826
rect 51490 9774 51492 9826
rect 51212 7028 51268 8372
rect 51212 6962 51268 6972
rect 50876 6626 50932 6636
rect 51436 6690 51492 9774
rect 51548 9716 51604 10332
rect 51660 10322 51716 10332
rect 51772 10052 51828 10062
rect 51884 10052 51940 10556
rect 51772 10050 51940 10052
rect 51772 9998 51774 10050
rect 51826 9998 51940 10050
rect 51772 9996 51940 9998
rect 51772 9986 51828 9996
rect 51548 9650 51604 9660
rect 51660 9602 51716 9614
rect 51660 9550 51662 9602
rect 51714 9550 51716 9602
rect 51660 8428 51716 9550
rect 51660 8372 51940 8428
rect 51884 8258 51940 8372
rect 51884 8206 51886 8258
rect 51938 8206 51940 8258
rect 51884 8194 51940 8206
rect 52108 8258 52164 12348
rect 52780 12338 52836 12348
rect 52892 23604 52948 23614
rect 52892 11844 52948 23548
rect 53564 23604 53620 102452
rect 53564 23538 53620 23548
rect 58156 21476 58212 21486
rect 57036 19124 57092 19134
rect 55804 14644 55860 14654
rect 52892 11778 52948 11788
rect 55132 12066 55188 12078
rect 55132 12014 55134 12066
rect 55186 12014 55188 12066
rect 54460 11508 54516 11518
rect 53788 11506 54516 11508
rect 53788 11454 54462 11506
rect 54514 11454 54516 11506
rect 53788 11452 54516 11454
rect 52780 11172 52836 11182
rect 53676 11172 53732 11182
rect 52444 10612 52500 10622
rect 52108 8206 52110 8258
rect 52162 8206 52164 8258
rect 52108 8194 52164 8206
rect 52220 10610 52500 10612
rect 52220 10558 52446 10610
rect 52498 10558 52500 10610
rect 52220 10556 52500 10558
rect 51436 6638 51438 6690
rect 51490 6638 51492 6690
rect 51324 6580 51380 6590
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 49980 5906 50036 5964
rect 49980 5854 49982 5906
rect 50034 5854 50036 5906
rect 49980 5842 50036 5854
rect 51212 5348 51268 5358
rect 49756 5236 49812 5246
rect 49756 5142 49812 5180
rect 49196 5010 49364 5012
rect 49196 4958 49198 5010
rect 49250 4958 49364 5010
rect 49196 4956 49364 4958
rect 49196 4946 49252 4956
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 49084 3614 49086 3666
rect 49138 3614 49140 3666
rect 49084 3602 49140 3614
rect 50876 4228 50932 4238
rect 49644 3444 49700 3454
rect 48748 3388 49140 3444
rect 47740 3350 47796 3388
rect 47516 1708 48020 1764
rect 47964 800 48020 1708
rect 49084 800 49140 3388
rect 49644 800 49700 3388
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50876 2996 50932 4172
rect 51212 3666 51268 5292
rect 51212 3614 51214 3666
rect 51266 3614 51268 3666
rect 51212 3602 51268 3614
rect 50764 2940 50932 2996
rect 50764 800 50820 2940
rect 51324 800 51380 6524
rect 51436 5236 51492 6638
rect 51436 5170 51492 5180
rect 51884 8036 51940 8046
rect 51884 5234 51940 7980
rect 52220 7924 52276 10556
rect 52444 10546 52500 10556
rect 52668 10612 52724 10622
rect 52332 10052 52388 10062
rect 52332 9826 52388 9996
rect 52668 10050 52724 10556
rect 52668 9998 52670 10050
rect 52722 9998 52724 10050
rect 52668 9986 52724 9998
rect 52332 9774 52334 9826
rect 52386 9774 52388 9826
rect 52332 9762 52388 9774
rect 52556 9602 52612 9614
rect 52556 9550 52558 9602
rect 52610 9550 52612 9602
rect 52444 8820 52500 8830
rect 52444 8258 52500 8764
rect 52444 8206 52446 8258
rect 52498 8206 52500 8258
rect 52444 8194 52500 8206
rect 52556 8260 52612 9550
rect 52780 8820 52836 11116
rect 53228 11170 53732 11172
rect 53228 11118 53678 11170
rect 53730 11118 53732 11170
rect 53228 11116 53732 11118
rect 53228 10722 53284 11116
rect 53676 11106 53732 11116
rect 53228 10670 53230 10722
rect 53282 10670 53284 10722
rect 53228 10658 53284 10670
rect 53564 10500 53620 10510
rect 53564 9154 53620 10444
rect 53676 9940 53732 9950
rect 53676 9846 53732 9884
rect 53564 9102 53566 9154
rect 53618 9102 53620 9154
rect 53564 9090 53620 9102
rect 52780 8754 52836 8764
rect 53340 8820 53396 8830
rect 52556 8194 52612 8204
rect 53340 8258 53396 8764
rect 53340 8206 53342 8258
rect 53394 8206 53396 8258
rect 53340 8194 53396 8206
rect 53788 8146 53844 11452
rect 54460 11442 54516 11452
rect 55020 11508 55076 11518
rect 55132 11508 55188 12014
rect 55020 11506 55188 11508
rect 55020 11454 55022 11506
rect 55074 11454 55188 11506
rect 55020 11452 55188 11454
rect 54012 11284 54068 11294
rect 54012 11282 54404 11284
rect 54012 11230 54014 11282
rect 54066 11230 54404 11282
rect 54012 11228 54404 11230
rect 54012 11218 54068 11228
rect 54348 10050 54404 11228
rect 54348 9998 54350 10050
rect 54402 9998 54404 10050
rect 54348 9986 54404 9998
rect 54684 10388 54740 10398
rect 54684 10050 54740 10332
rect 54684 9998 54686 10050
rect 54738 9998 54740 10050
rect 54684 9986 54740 9998
rect 53788 8094 53790 8146
rect 53842 8094 53844 8146
rect 52332 8036 52388 8046
rect 52332 7942 52388 7980
rect 53564 8034 53620 8046
rect 53564 7982 53566 8034
rect 53618 7982 53620 8034
rect 51884 5182 51886 5234
rect 51938 5182 51940 5234
rect 51884 5170 51940 5182
rect 52108 6804 52164 6814
rect 51996 4676 52052 4686
rect 51996 4450 52052 4620
rect 51996 4398 51998 4450
rect 52050 4398 52052 4450
rect 51996 4340 52052 4398
rect 51996 3554 52052 4284
rect 51996 3502 51998 3554
rect 52050 3502 52052 3554
rect 51996 3490 52052 3502
rect 52108 2884 52164 6748
rect 52220 6692 52276 7868
rect 52220 6020 52276 6636
rect 53452 6692 53508 6702
rect 53452 6598 53508 6636
rect 52332 6580 52388 6590
rect 52332 6486 52388 6524
rect 52220 6018 52612 6020
rect 52220 5966 52222 6018
rect 52274 5966 52612 6018
rect 52220 5964 52612 5966
rect 52220 5954 52276 5964
rect 52108 2818 52164 2828
rect 52444 5684 52500 5694
rect 52444 800 52500 5628
rect 52556 5124 52612 5964
rect 53564 5348 53620 7982
rect 53788 6804 53844 8094
rect 53788 6738 53844 6748
rect 53900 9940 53956 9950
rect 53900 9044 53956 9884
rect 55020 9940 55076 11452
rect 55468 11172 55524 11182
rect 55356 10500 55412 10510
rect 55020 9268 55076 9884
rect 55244 10498 55412 10500
rect 55244 10446 55358 10498
rect 55410 10446 55412 10498
rect 55244 10444 55412 10446
rect 55244 9716 55300 10444
rect 55356 10434 55412 10444
rect 55468 10276 55524 11116
rect 55020 9202 55076 9212
rect 55132 9714 55300 9716
rect 55132 9662 55246 9714
rect 55298 9662 55300 9714
rect 55132 9660 55300 9662
rect 53900 7474 53956 8988
rect 54796 9044 54852 9054
rect 54012 8260 54068 8270
rect 54012 8166 54068 8204
rect 54796 8258 54852 8988
rect 55132 8428 55188 9660
rect 55244 9650 55300 9660
rect 55356 10220 55524 10276
rect 55580 11170 55636 11182
rect 55580 11118 55582 11170
rect 55634 11118 55636 11170
rect 54796 8206 54798 8258
rect 54850 8206 54852 8258
rect 53900 7422 53902 7474
rect 53954 7422 53956 7474
rect 53564 5282 53620 5292
rect 52556 4992 52612 5068
rect 53788 5124 53844 5134
rect 53788 5030 53844 5068
rect 53900 4338 53956 7422
rect 54236 8036 54292 8046
rect 54236 6690 54292 7980
rect 54236 6638 54238 6690
rect 54290 6638 54292 6690
rect 54236 6626 54292 6638
rect 54796 6244 54852 8206
rect 54796 6178 54852 6188
rect 54908 8372 55188 8428
rect 55244 9156 55300 9166
rect 54908 6020 54964 8372
rect 55244 8370 55300 9100
rect 55244 8318 55246 8370
rect 55298 8318 55300 8370
rect 55244 8306 55300 8318
rect 55356 9154 55412 10220
rect 55356 9102 55358 9154
rect 55410 9102 55412 9154
rect 55356 7700 55412 9102
rect 55244 7644 55412 7700
rect 55468 9826 55524 9838
rect 55468 9774 55470 9826
rect 55522 9774 55524 9826
rect 55468 9156 55524 9774
rect 55244 6468 55300 7644
rect 55356 7476 55412 7486
rect 55356 7382 55412 7420
rect 55244 6402 55300 6412
rect 54124 5964 54964 6020
rect 53900 4286 53902 4338
rect 53954 4286 53956 4338
rect 53900 4274 53956 4286
rect 54012 5012 54068 5022
rect 53116 3668 53172 3678
rect 53004 3666 53172 3668
rect 53004 3614 53118 3666
rect 53170 3614 53172 3666
rect 53004 3612 53172 3614
rect 53004 800 53060 3612
rect 53116 3602 53172 3612
rect 54012 3332 54068 4956
rect 54124 3554 54180 5964
rect 55468 5906 55524 9100
rect 55580 7476 55636 11118
rect 55692 9604 55748 9614
rect 55692 9266 55748 9548
rect 55692 9214 55694 9266
rect 55746 9214 55748 9266
rect 55692 9044 55748 9214
rect 55692 8978 55748 8988
rect 55692 7700 55748 7710
rect 55804 7700 55860 14588
rect 56588 13972 56644 13982
rect 56252 12516 56308 12526
rect 56140 11620 56196 11630
rect 56028 11172 56084 11182
rect 56028 11078 56084 11116
rect 56028 10836 56084 10846
rect 56140 10836 56196 11564
rect 56028 10834 56196 10836
rect 56028 10782 56030 10834
rect 56082 10782 56196 10834
rect 56028 10780 56196 10782
rect 55916 10612 55972 10622
rect 55916 8428 55972 10556
rect 56028 10388 56084 10780
rect 56028 10322 56084 10332
rect 56140 10500 56196 10510
rect 56140 9826 56196 10444
rect 56140 9774 56142 9826
rect 56194 9774 56196 9826
rect 56140 9762 56196 9774
rect 56140 9044 56196 9054
rect 56140 8950 56196 8988
rect 56252 8428 56308 12460
rect 56364 11170 56420 11182
rect 56364 11118 56366 11170
rect 56418 11118 56420 11170
rect 56364 9604 56420 11118
rect 56476 10500 56532 10510
rect 56476 10406 56532 10444
rect 56364 9538 56420 9548
rect 55916 8372 56084 8428
rect 55916 8036 55972 8046
rect 55916 7942 55972 7980
rect 55692 7698 55860 7700
rect 55692 7646 55694 7698
rect 55746 7646 55860 7698
rect 55692 7644 55860 7646
rect 55692 7634 55748 7644
rect 56028 7586 56084 8372
rect 56028 7534 56030 7586
rect 56082 7534 56084 7586
rect 56028 7522 56084 7534
rect 56140 8372 56308 8428
rect 55580 7410 55636 7420
rect 55804 7476 55860 7486
rect 55468 5854 55470 5906
rect 55522 5854 55524 5906
rect 55468 5842 55524 5854
rect 55692 6020 55748 6030
rect 54572 5236 54628 5246
rect 54572 5142 54628 5180
rect 54124 3502 54126 3554
rect 54178 3502 54180 3554
rect 54124 3490 54180 3502
rect 54684 4228 54740 4238
rect 54012 3276 54180 3332
rect 54124 800 54180 3276
rect 54684 800 54740 4172
rect 55580 4228 55636 4238
rect 55580 4134 55636 4172
rect 55692 3554 55748 5964
rect 55692 3502 55694 3554
rect 55746 3502 55748 3554
rect 55692 3490 55748 3502
rect 55020 3444 55076 3454
rect 55020 3350 55076 3388
rect 55804 800 55860 7420
rect 56140 5908 56196 8372
rect 56252 8148 56308 8158
rect 56252 8146 56532 8148
rect 56252 8094 56254 8146
rect 56306 8094 56532 8146
rect 56252 8092 56532 8094
rect 56252 8082 56308 8092
rect 56252 7588 56308 7598
rect 56252 7586 56420 7588
rect 56252 7534 56254 7586
rect 56306 7534 56420 7586
rect 56252 7532 56420 7534
rect 56252 7522 56308 7532
rect 56364 7474 56420 7532
rect 56364 7422 56366 7474
rect 56418 7422 56420 7474
rect 56364 7410 56420 7422
rect 56364 6802 56420 6814
rect 56364 6750 56366 6802
rect 56418 6750 56420 6802
rect 56364 6020 56420 6750
rect 56476 6132 56532 8092
rect 56588 6580 56644 13916
rect 57036 12516 57092 19068
rect 57036 12450 57092 12460
rect 57708 15988 57764 15998
rect 57372 12292 57428 12302
rect 57372 12198 57428 12236
rect 57260 11954 57316 11966
rect 57260 11902 57262 11954
rect 57314 11902 57316 11954
rect 57148 11618 57204 11630
rect 57148 11566 57150 11618
rect 57202 11566 57204 11618
rect 56812 11170 56868 11182
rect 56812 11118 56814 11170
rect 56866 11118 56868 11170
rect 56812 10612 56868 11118
rect 56812 10546 56868 10556
rect 56924 10724 56980 10734
rect 56924 9938 56980 10668
rect 56924 9886 56926 9938
rect 56978 9886 56980 9938
rect 56924 9874 56980 9886
rect 56700 9044 56756 9054
rect 56700 8950 56756 8988
rect 57036 8034 57092 8046
rect 57036 7982 57038 8034
rect 57090 7982 57092 8034
rect 57036 7700 57092 7982
rect 57036 7634 57092 7644
rect 56700 7476 56756 7486
rect 56700 7474 56868 7476
rect 56700 7422 56702 7474
rect 56754 7422 56868 7474
rect 56700 7420 56868 7422
rect 56700 7410 56756 7420
rect 56588 6514 56644 6524
rect 56700 7250 56756 7262
rect 56700 7198 56702 7250
rect 56754 7198 56756 7250
rect 56588 6132 56644 6142
rect 56476 6130 56644 6132
rect 56476 6078 56590 6130
rect 56642 6078 56644 6130
rect 56476 6076 56644 6078
rect 56588 6066 56644 6076
rect 56364 5954 56420 5964
rect 56700 6020 56756 7198
rect 56700 5954 56756 5964
rect 56252 5908 56308 5918
rect 56140 5906 56308 5908
rect 56140 5854 56254 5906
rect 56306 5854 56308 5906
rect 56140 5852 56308 5854
rect 56252 5842 56308 5852
rect 56700 5236 56756 5246
rect 56812 5236 56868 7420
rect 57148 7140 57204 11566
rect 57148 7074 57204 7084
rect 56700 5234 56868 5236
rect 56700 5182 56702 5234
rect 56754 5182 56868 5234
rect 56700 5180 56868 5182
rect 57148 6692 57204 6702
rect 56588 4340 56644 4350
rect 56700 4340 56756 5180
rect 56588 4338 56756 4340
rect 56588 4286 56590 4338
rect 56642 4286 56756 4338
rect 56588 4284 56756 4286
rect 57036 5124 57092 5134
rect 57036 4788 57092 5068
rect 57148 5012 57204 6636
rect 57260 5124 57316 11902
rect 57484 11172 57540 11182
rect 57484 11170 57652 11172
rect 57484 11118 57486 11170
rect 57538 11118 57652 11170
rect 57484 11116 57652 11118
rect 57484 11106 57540 11116
rect 57484 10724 57540 10734
rect 57484 10630 57540 10668
rect 57484 8146 57540 8158
rect 57484 8094 57486 8146
rect 57538 8094 57540 8146
rect 57484 7700 57540 8094
rect 57484 7634 57540 7644
rect 57596 6580 57652 11116
rect 57708 8148 57764 15932
rect 57932 12516 57988 12526
rect 57932 12402 57988 12460
rect 57932 12350 57934 12402
rect 57986 12350 57988 12402
rect 57932 12338 57988 12350
rect 57932 11618 57988 11630
rect 57932 11566 57934 11618
rect 57986 11566 57988 11618
rect 57932 11506 57988 11566
rect 57932 11454 57934 11506
rect 57986 11454 57988 11506
rect 57932 11442 57988 11454
rect 57820 10610 57876 10622
rect 57820 10558 57822 10610
rect 57874 10558 57876 10610
rect 57820 9268 57876 10558
rect 58044 10386 58100 10398
rect 58044 10334 58046 10386
rect 58098 10334 58100 10386
rect 57932 9268 57988 9278
rect 57820 9266 57988 9268
rect 57820 9214 57934 9266
rect 57986 9214 57988 9266
rect 57820 9212 57988 9214
rect 57932 9202 57988 9212
rect 57820 8148 57876 8158
rect 57708 8146 57876 8148
rect 57708 8094 57822 8146
rect 57874 8094 57876 8146
rect 57708 8092 57876 8094
rect 57820 8082 57876 8092
rect 57820 7476 57876 7486
rect 58044 7476 58100 10334
rect 57820 7474 58100 7476
rect 57820 7422 57822 7474
rect 57874 7422 58100 7474
rect 57820 7420 58100 7422
rect 57708 6580 57764 6590
rect 57596 6578 57764 6580
rect 57596 6526 57710 6578
rect 57762 6526 57764 6578
rect 57596 6524 57764 6526
rect 57484 6020 57540 6030
rect 57484 5926 57540 5964
rect 57260 5068 57428 5124
rect 57148 4946 57204 4956
rect 57260 4898 57316 4910
rect 57260 4846 57262 4898
rect 57314 4846 57316 4898
rect 57260 4788 57316 4846
rect 57036 4732 57316 4788
rect 56588 4274 56644 4284
rect 56364 3444 56420 3454
rect 56364 800 56420 3388
rect 57036 2772 57092 4732
rect 57372 4340 57428 5068
rect 57484 4340 57540 4350
rect 57372 4284 57484 4340
rect 57484 4246 57540 4284
rect 57596 4116 57652 6524
rect 57708 6514 57764 6524
rect 57708 6020 57764 6030
rect 57708 5926 57764 5964
rect 57708 5124 57764 5134
rect 57820 5124 57876 7420
rect 57932 7140 57988 7150
rect 57932 6020 57988 7084
rect 58044 6580 58100 6590
rect 58044 6486 58100 6524
rect 58044 6020 58100 6030
rect 57932 6018 58100 6020
rect 57932 5966 58046 6018
rect 58098 5966 58100 6018
rect 57932 5964 58100 5966
rect 58044 5954 58100 5964
rect 57932 5794 57988 5806
rect 57932 5742 57934 5794
rect 57986 5742 57988 5794
rect 57932 5236 57988 5742
rect 57932 5170 57988 5180
rect 57708 5122 57876 5124
rect 57708 5070 57710 5122
rect 57762 5070 57876 5122
rect 57708 5068 57876 5070
rect 57708 4676 57764 5068
rect 57708 4610 57764 4620
rect 57820 4564 57876 4574
rect 58156 4564 58212 21420
rect 62860 19460 62916 116174
rect 64092 116004 64148 119200
rect 65660 116676 65716 119200
rect 68796 117572 68852 119200
rect 68796 117516 69300 117572
rect 65916 116844 66180 116854
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 65916 116778 66180 116788
rect 65660 116620 66164 116676
rect 66108 116562 66164 116620
rect 66108 116510 66110 116562
rect 66162 116510 66164 116562
rect 66108 116498 66164 116510
rect 69244 116562 69300 117516
rect 69244 116510 69246 116562
rect 69298 116510 69300 116562
rect 69244 116498 69300 116510
rect 70364 116564 70420 119200
rect 70588 116564 70644 116574
rect 70364 116562 70644 116564
rect 70364 116510 70590 116562
rect 70642 116510 70644 116562
rect 70364 116508 70644 116510
rect 70588 116498 70644 116508
rect 73052 116564 73108 116574
rect 67116 116450 67172 116462
rect 67116 116398 67118 116450
rect 67170 116398 67172 116450
rect 67116 116228 67172 116398
rect 68796 116450 68852 116462
rect 68796 116398 68798 116450
rect 68850 116398 68852 116450
rect 67116 116162 67172 116172
rect 67564 116228 67620 116238
rect 67564 116134 67620 116172
rect 64092 115948 64260 116004
rect 64092 115778 64148 115790
rect 64092 115726 64094 115778
rect 64146 115726 64148 115778
rect 63756 115666 63812 115678
rect 63756 115614 63758 115666
rect 63810 115614 63812 115666
rect 63196 115556 63252 115566
rect 63196 115462 63252 115500
rect 63756 115556 63812 115614
rect 63756 115490 63812 115500
rect 64092 114884 64148 115726
rect 64204 115108 64260 115948
rect 68796 115890 68852 116398
rect 71372 116450 71428 116462
rect 71372 116398 71374 116450
rect 71426 116398 71428 116450
rect 68796 115838 68798 115890
rect 68850 115838 68852 115890
rect 68796 115826 68852 115838
rect 69916 116228 69972 116238
rect 68572 115666 68628 115678
rect 68572 115614 68574 115666
rect 68626 115614 68628 115666
rect 67900 115556 67956 115566
rect 67900 115462 67956 115500
rect 68572 115556 68628 115614
rect 68572 115490 68628 115500
rect 65916 115276 66180 115286
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 65916 115210 66180 115220
rect 64204 115042 64260 115052
rect 64988 115108 65044 115118
rect 64988 114994 65044 115052
rect 64988 114942 64990 114994
rect 65042 114942 65044 114994
rect 64988 114930 65044 114942
rect 64316 114884 64372 114894
rect 64092 114882 64372 114884
rect 64092 114830 64318 114882
rect 64370 114830 64372 114882
rect 64092 114828 64372 114830
rect 64316 114818 64372 114828
rect 65916 113708 66180 113718
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 65916 113642 66180 113652
rect 65916 112140 66180 112150
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 65916 112074 66180 112084
rect 65916 110572 66180 110582
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 65916 110506 66180 110516
rect 65916 109004 66180 109014
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 65916 108938 66180 108948
rect 65916 107436 66180 107446
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 65916 107370 66180 107380
rect 65916 105868 66180 105878
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 65916 105802 66180 105812
rect 65916 104300 66180 104310
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 65916 104234 66180 104244
rect 65916 102732 66180 102742
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 65916 102666 66180 102676
rect 65916 101164 66180 101174
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 65916 101098 66180 101108
rect 65916 99596 66180 99606
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 65916 99530 66180 99540
rect 65916 98028 66180 98038
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 65916 97962 66180 97972
rect 65916 96460 66180 96470
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 65916 96394 66180 96404
rect 65916 94892 66180 94902
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 65916 94826 66180 94836
rect 65916 93324 66180 93334
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 65916 93258 66180 93268
rect 65916 91756 66180 91766
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 65916 91690 66180 91700
rect 65916 90188 66180 90198
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 65916 90122 66180 90132
rect 65916 88620 66180 88630
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 65916 88554 66180 88564
rect 65916 87052 66180 87062
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 65916 86986 66180 86996
rect 65916 85484 66180 85494
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 65916 85418 66180 85428
rect 65916 83916 66180 83926
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 65916 83850 66180 83860
rect 65916 82348 66180 82358
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 65916 82282 66180 82292
rect 65916 80780 66180 80790
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 65916 80714 66180 80724
rect 65916 79212 66180 79222
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 65916 79146 66180 79156
rect 65916 77644 66180 77654
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 65916 77578 66180 77588
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 67900 27412 67956 27422
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 62860 19394 62916 19404
rect 65548 24164 65604 24174
rect 63756 19348 63812 19358
rect 58492 19012 58548 19022
rect 58380 12066 58436 12078
rect 58380 12014 58382 12066
rect 58434 12014 58436 12066
rect 58380 11954 58436 12014
rect 58380 11902 58382 11954
rect 58434 11902 58436 11954
rect 58380 11890 58436 11902
rect 58380 11508 58436 11518
rect 58492 11508 58548 18956
rect 62188 17444 62244 17454
rect 58940 16212 58996 16222
rect 58380 11506 58548 11508
rect 58380 11454 58382 11506
rect 58434 11454 58548 11506
rect 58380 11452 58548 11454
rect 58604 12292 58660 12302
rect 58268 10498 58324 10510
rect 58268 10446 58270 10498
rect 58322 10446 58324 10498
rect 58268 10386 58324 10446
rect 58268 10334 58270 10386
rect 58322 10334 58324 10386
rect 58268 10322 58324 10334
rect 58268 8932 58324 8942
rect 58268 8838 58324 8876
rect 58380 8428 58436 11452
rect 58268 8372 58436 8428
rect 58492 9156 58548 9166
rect 58268 6020 58324 8372
rect 58380 8036 58436 8046
rect 58380 7942 58436 7980
rect 58492 6020 58548 9100
rect 58604 9154 58660 12236
rect 58716 11170 58772 11182
rect 58716 11118 58718 11170
rect 58770 11118 58772 11170
rect 58716 10386 58772 11118
rect 58716 10334 58718 10386
rect 58770 10334 58772 10386
rect 58716 10322 58772 10334
rect 58828 10498 58884 10510
rect 58828 10446 58830 10498
rect 58882 10446 58884 10498
rect 58828 9380 58884 10446
rect 58604 9102 58606 9154
rect 58658 9102 58660 9154
rect 58604 9044 58660 9102
rect 58604 8978 58660 8988
rect 58716 9324 58884 9380
rect 58716 8932 58772 9324
rect 58828 9156 58884 9166
rect 58828 9062 58884 9100
rect 58716 8876 58884 8932
rect 58716 8036 58772 8046
rect 58604 7362 58660 7374
rect 58604 7310 58606 7362
rect 58658 7310 58660 7362
rect 58604 6356 58660 7310
rect 58716 6580 58772 7980
rect 58828 6692 58884 8876
rect 58940 8036 58996 16156
rect 61740 14756 61796 14766
rect 60508 14532 60564 14542
rect 59612 12292 59668 12302
rect 59612 12198 59668 12236
rect 59164 12068 59220 12078
rect 59164 11732 59220 12012
rect 60284 11956 60340 11966
rect 60172 11954 60340 11956
rect 60172 11902 60286 11954
rect 60338 11902 60340 11954
rect 60172 11900 60340 11902
rect 59164 11676 59556 11732
rect 59388 11508 59444 11518
rect 59052 9938 59108 9950
rect 59052 9886 59054 9938
rect 59106 9886 59108 9938
rect 59052 9156 59108 9886
rect 59052 9090 59108 9100
rect 59276 8484 59332 8494
rect 59276 8260 59332 8428
rect 59388 8428 59444 11452
rect 59500 10498 59556 11676
rect 59948 11508 60004 11518
rect 59948 11414 60004 11452
rect 59500 10446 59502 10498
rect 59554 10446 59556 10498
rect 59500 10388 59556 10446
rect 59500 10332 60004 10388
rect 59612 9604 59668 9614
rect 59500 9602 59668 9604
rect 59500 9550 59614 9602
rect 59666 9550 59668 9602
rect 59500 9548 59668 9550
rect 59500 8596 59556 9548
rect 59612 9538 59668 9548
rect 59948 9604 60004 10332
rect 60172 9826 60228 11900
rect 60284 11890 60340 11900
rect 60508 11508 60564 14476
rect 61516 13636 61572 13646
rect 60844 12292 60900 12302
rect 60844 12198 60900 12236
rect 61180 12290 61236 12302
rect 61180 12238 61182 12290
rect 61234 12238 61236 12290
rect 61180 12068 61236 12238
rect 61180 12002 61236 12012
rect 60620 11956 60676 11966
rect 60620 11862 60676 11900
rect 60508 11442 60564 11452
rect 60172 9774 60174 9826
rect 60226 9774 60228 9826
rect 60172 9762 60228 9774
rect 60284 11170 60340 11182
rect 61292 11172 61348 11182
rect 60284 11118 60286 11170
rect 60338 11118 60340 11170
rect 60284 9604 60340 11118
rect 61068 11170 61348 11172
rect 61068 11118 61294 11170
rect 61346 11118 61348 11170
rect 61068 11116 61348 11118
rect 60508 10612 60564 10622
rect 60508 9714 60564 10556
rect 60508 9662 60510 9714
rect 60562 9662 60564 9714
rect 60508 9650 60564 9662
rect 59948 9548 60340 9604
rect 59612 9156 59668 9166
rect 59612 9062 59668 9100
rect 59500 8540 59668 8596
rect 59612 8428 59668 8540
rect 59724 8482 59780 8494
rect 59724 8430 59726 8482
rect 59778 8430 59780 8482
rect 59724 8428 59780 8430
rect 59948 8428 60004 9548
rect 60620 9044 60676 9054
rect 60620 8950 60676 8988
rect 59388 8372 59556 8428
rect 59612 8372 59780 8428
rect 59276 8166 59332 8204
rect 58940 7942 58996 7980
rect 59164 7700 59220 7710
rect 58828 6636 58996 6692
rect 58716 6524 58884 6580
rect 58828 6466 58884 6524
rect 58828 6414 58830 6466
rect 58882 6414 58884 6466
rect 58828 6402 58884 6414
rect 58604 6290 58660 6300
rect 58268 5954 58324 5964
rect 58380 5964 58548 6020
rect 57820 4562 58212 4564
rect 57820 4510 57822 4562
rect 57874 4510 58212 4562
rect 57820 4508 58212 4510
rect 57820 4498 57876 4508
rect 58380 4452 58436 5964
rect 58940 5906 58996 6636
rect 58940 5854 58942 5906
rect 58994 5854 58996 5906
rect 58604 5794 58660 5806
rect 58604 5742 58606 5794
rect 58658 5742 58660 5794
rect 58604 5684 58660 5742
rect 58604 5618 58660 5628
rect 58492 5236 58548 5246
rect 58492 5142 58548 5180
rect 58940 4564 58996 5854
rect 58940 4498 58996 4508
rect 57484 4060 57652 4116
rect 57932 4396 58436 4452
rect 57148 3444 57204 3454
rect 57148 3350 57204 3388
rect 57036 2706 57092 2716
rect 57484 800 57540 4060
rect 57932 3554 57988 4396
rect 57932 3502 57934 3554
rect 57986 3502 57988 3554
rect 57932 3490 57988 3502
rect 58380 4226 58436 4238
rect 58380 4174 58382 4226
rect 58434 4174 58436 4226
rect 58044 3444 58100 3454
rect 58044 800 58100 3388
rect 58380 3332 58436 4174
rect 58940 3444 58996 3454
rect 58940 3350 58996 3388
rect 58380 2660 58436 3276
rect 58380 2594 58436 2604
rect 59164 800 59220 7644
rect 59388 6580 59444 6590
rect 59388 6486 59444 6524
rect 59388 6132 59444 6142
rect 59500 6132 59556 8372
rect 59724 8034 59780 8372
rect 59724 7982 59726 8034
rect 59778 7982 59780 8034
rect 59724 7140 59780 7982
rect 59724 6692 59780 7084
rect 59724 6626 59780 6636
rect 59836 8372 60004 8428
rect 60060 8482 60116 8494
rect 60060 8430 60062 8482
rect 60114 8430 60116 8482
rect 60060 8428 60116 8430
rect 60060 8372 60228 8428
rect 59388 6130 59556 6132
rect 59388 6078 59390 6130
rect 59442 6078 59556 6130
rect 59388 6076 59556 6078
rect 59724 6466 59780 6478
rect 59724 6414 59726 6466
rect 59778 6414 59780 6466
rect 59388 6066 59444 6076
rect 59612 5908 59668 5918
rect 59612 5814 59668 5852
rect 59500 5794 59556 5806
rect 59500 5742 59502 5794
rect 59554 5742 59556 5794
rect 59500 5236 59556 5742
rect 59500 5170 59556 5180
rect 59724 4452 59780 6414
rect 59724 4386 59780 4396
rect 59836 3554 59892 8372
rect 60172 8370 60228 8372
rect 60172 8318 60174 8370
rect 60226 8318 60228 8370
rect 60172 8306 60228 8318
rect 60732 8034 60788 8046
rect 60732 7982 60734 8034
rect 60786 7982 60788 8034
rect 60732 7588 60788 7982
rect 60732 7522 60788 7532
rect 60956 7588 61012 7598
rect 60732 7364 60788 7374
rect 60732 7362 60900 7364
rect 60732 7310 60734 7362
rect 60786 7310 60900 7362
rect 60732 7308 60900 7310
rect 60732 7298 60788 7308
rect 60620 6578 60676 6590
rect 60620 6526 60622 6578
rect 60674 6526 60676 6578
rect 60396 6468 60452 6478
rect 60396 6374 60452 6412
rect 60508 6466 60564 6478
rect 60508 6414 60510 6466
rect 60562 6414 60564 6466
rect 60396 6132 60452 6142
rect 60396 5906 60452 6076
rect 60508 6020 60564 6414
rect 60620 6244 60676 6526
rect 60620 6178 60676 6188
rect 60844 6468 60900 7308
rect 60508 5954 60564 5964
rect 60732 6018 60788 6030
rect 60732 5966 60734 6018
rect 60786 5966 60788 6018
rect 60396 5854 60398 5906
rect 60450 5854 60452 5906
rect 60396 5124 60452 5854
rect 60620 5234 60676 5246
rect 60620 5182 60622 5234
rect 60674 5182 60676 5234
rect 60396 5068 60564 5124
rect 60508 4788 60564 5068
rect 60620 5012 60676 5182
rect 60620 4946 60676 4956
rect 60508 4732 60676 4788
rect 60508 4452 60564 4462
rect 60508 4358 60564 4396
rect 59836 3502 59838 3554
rect 59890 3502 59892 3554
rect 59836 3490 59892 3502
rect 59724 3444 59780 3454
rect 59724 800 59780 3388
rect 60620 1316 60676 4732
rect 60732 1540 60788 5966
rect 60844 3554 60900 6412
rect 60956 4564 61012 7532
rect 61068 6132 61124 11116
rect 61292 11106 61348 11116
rect 61516 10836 61572 13580
rect 61068 6066 61124 6076
rect 61180 9044 61236 9054
rect 60956 4498 61012 4508
rect 61180 4338 61236 8988
rect 61292 8930 61348 8942
rect 61292 8878 61294 8930
rect 61346 8878 61348 8930
rect 61292 7700 61348 8878
rect 61516 8428 61572 10780
rect 61628 10612 61684 10650
rect 61628 10546 61684 10556
rect 61740 10276 61796 14700
rect 61964 12066 62020 12078
rect 61964 12014 61966 12066
rect 62018 12014 62020 12066
rect 61964 11956 62020 12014
rect 61964 11890 62020 11900
rect 62188 11396 62244 17388
rect 62076 11340 62244 11396
rect 63420 16324 63476 16334
rect 61628 10220 61796 10276
rect 61852 11170 61908 11182
rect 61852 11118 61854 11170
rect 61906 11118 61908 11170
rect 61628 9156 61684 10220
rect 61740 10050 61796 10062
rect 61740 9998 61742 10050
rect 61794 9998 61796 10050
rect 61740 9938 61796 9998
rect 61740 9886 61742 9938
rect 61794 9886 61796 9938
rect 61740 9874 61796 9886
rect 61628 9090 61684 9100
rect 61852 8428 61908 11118
rect 62076 10500 62132 11340
rect 62188 11170 62244 11182
rect 62188 11118 62190 11170
rect 62242 11118 62244 11170
rect 62188 10612 62244 11118
rect 62636 11170 62692 11182
rect 62636 11118 62638 11170
rect 62690 11118 62692 11170
rect 62636 11060 62692 11118
rect 62636 10994 62692 11004
rect 63196 11172 63252 11182
rect 62300 10612 62356 10622
rect 62188 10610 62356 10612
rect 62188 10558 62302 10610
rect 62354 10558 62356 10610
rect 62188 10556 62356 10558
rect 62300 10500 62356 10556
rect 62860 10500 62916 10510
rect 62076 10444 62244 10500
rect 62076 10050 62132 10062
rect 62076 9998 62078 10050
rect 62130 9998 62132 10050
rect 61516 8372 61796 8428
rect 61852 8372 62020 8428
rect 61404 8260 61460 8270
rect 61404 8166 61460 8204
rect 61292 7634 61348 7644
rect 61516 8036 61572 8046
rect 61404 7364 61460 7374
rect 61292 6020 61348 6030
rect 61292 5926 61348 5964
rect 61404 4900 61460 7308
rect 61516 6018 61572 7980
rect 61740 7698 61796 8372
rect 61740 7646 61742 7698
rect 61794 7646 61796 7698
rect 61740 7634 61796 7646
rect 61852 6692 61908 6702
rect 61740 6468 61796 6478
rect 61740 6374 61796 6412
rect 61628 6356 61684 6366
rect 61628 6130 61684 6300
rect 61628 6078 61630 6130
rect 61682 6078 61684 6130
rect 61628 6066 61684 6078
rect 61516 5966 61518 6018
rect 61570 5966 61572 6018
rect 61516 5954 61572 5966
rect 61852 6018 61908 6636
rect 61852 5966 61854 6018
rect 61906 5966 61908 6018
rect 61852 5954 61908 5966
rect 61964 5796 62020 8372
rect 61740 5740 62020 5796
rect 61404 4834 61460 4844
rect 61516 5012 61572 5022
rect 61740 5012 61796 5740
rect 61852 5124 61908 5134
rect 61852 5030 61908 5068
rect 61516 5010 61796 5012
rect 61516 4958 61518 5010
rect 61570 4958 61796 5010
rect 61516 4956 61796 4958
rect 61180 4286 61182 4338
rect 61234 4286 61236 4338
rect 61180 4274 61236 4286
rect 60844 3502 60846 3554
rect 60898 3502 60900 3554
rect 60844 3490 60900 3502
rect 61404 3666 61460 3678
rect 61404 3614 61406 3666
rect 61458 3614 61460 3666
rect 60732 1474 60788 1484
rect 60620 1260 60900 1316
rect 60844 800 60900 1260
rect 61404 800 61460 3614
rect 61516 3332 61572 4956
rect 61852 4564 61908 4574
rect 61852 4470 61908 4508
rect 62076 4452 62132 9998
rect 62188 9938 62244 10444
rect 62188 9886 62190 9938
rect 62242 9886 62244 9938
rect 62188 8820 62244 9886
rect 62300 10498 62916 10500
rect 62300 10446 62862 10498
rect 62914 10446 62916 10498
rect 62300 10444 62916 10446
rect 62300 9940 62356 10444
rect 62860 10434 62916 10444
rect 62300 9044 62356 9884
rect 62636 10164 62692 10174
rect 62300 8978 62356 8988
rect 62524 9604 62580 9614
rect 62524 9044 62580 9548
rect 62524 8978 62580 8988
rect 62188 8764 62580 8820
rect 62188 8484 62244 8494
rect 62188 6690 62244 8428
rect 62412 7700 62468 7710
rect 62412 7606 62468 7644
rect 62188 6638 62190 6690
rect 62242 6638 62244 6690
rect 62188 6626 62244 6638
rect 62300 7474 62356 7486
rect 62300 7422 62302 7474
rect 62354 7422 62356 7474
rect 62300 6692 62356 7422
rect 62524 7474 62580 8764
rect 62524 7422 62526 7474
rect 62578 7422 62580 7474
rect 62524 7410 62580 7422
rect 62636 6804 62692 10108
rect 63196 10164 63252 11116
rect 63420 10836 63476 16268
rect 63756 12964 63812 19292
rect 63756 12908 64260 12964
rect 63756 12292 63812 12302
rect 63756 12198 63812 12236
rect 63756 11508 63812 11518
rect 63868 11508 63924 12908
rect 64204 12402 64260 12908
rect 64204 12350 64206 12402
rect 64258 12350 64260 12402
rect 64204 12338 64260 12350
rect 63812 11452 63924 11508
rect 64540 12292 64596 12302
rect 63756 11376 63812 11452
rect 63980 11396 64036 11406
rect 63420 10834 63700 10836
rect 63420 10782 63422 10834
rect 63474 10782 63700 10834
rect 63420 10780 63700 10782
rect 63420 10770 63476 10780
rect 63196 10098 63252 10108
rect 63420 9940 63476 9950
rect 63420 9846 63476 9884
rect 62972 9604 63028 9614
rect 62972 9510 63028 9548
rect 63420 9044 63476 9054
rect 62860 8932 62916 8942
rect 62860 7586 62916 8876
rect 63420 8930 63476 8988
rect 63420 8878 63422 8930
rect 63474 8878 63476 8930
rect 63420 8428 63476 8878
rect 62860 7534 62862 7586
rect 62914 7534 62916 7586
rect 62860 7522 62916 7534
rect 63308 8372 63476 8428
rect 62300 6626 62356 6636
rect 62524 6748 62692 6804
rect 62972 7028 63028 7038
rect 62972 6802 63028 6972
rect 62972 6750 62974 6802
rect 63026 6750 63028 6802
rect 62524 5906 62580 6748
rect 62972 6738 63028 6750
rect 62524 5854 62526 5906
rect 62578 5854 62580 5906
rect 62300 5348 62356 5358
rect 62300 5254 62356 5292
rect 62524 5012 62580 5854
rect 62636 6580 62692 6590
rect 62636 5346 62692 6524
rect 62860 6356 62916 6366
rect 62860 6130 62916 6300
rect 62860 6078 62862 6130
rect 62914 6078 62916 6130
rect 62636 5294 62638 5346
rect 62690 5294 62692 5346
rect 62636 5282 62692 5294
rect 62748 5348 62804 5358
rect 62524 4946 62580 4956
rect 62076 4386 62132 4396
rect 62300 4676 62356 4686
rect 62300 4450 62356 4620
rect 62636 4564 62692 4574
rect 62748 4564 62804 5292
rect 62860 5124 62916 6078
rect 62860 5058 62916 5068
rect 62636 4562 62804 4564
rect 62636 4510 62638 4562
rect 62690 4510 62804 4562
rect 62636 4508 62804 4510
rect 63196 4900 63252 4910
rect 62636 4498 62692 4508
rect 62300 4398 62302 4450
rect 62354 4398 62356 4450
rect 62300 4386 62356 4398
rect 63196 4450 63252 4844
rect 63196 4398 63198 4450
rect 63250 4398 63252 4450
rect 63196 4386 63252 4398
rect 61516 3266 61572 3276
rect 62524 4340 62580 4350
rect 62524 800 62580 4284
rect 63084 3666 63140 3678
rect 63084 3614 63086 3666
rect 63138 3614 63140 3666
rect 63084 800 63140 3614
rect 63308 3556 63364 8372
rect 63420 7474 63476 7486
rect 63420 7422 63422 7474
rect 63474 7422 63476 7474
rect 63420 6692 63476 7422
rect 63644 7474 63700 10780
rect 63980 10612 64036 11340
rect 63756 10498 63812 10510
rect 63756 10446 63758 10498
rect 63810 10446 63812 10498
rect 63756 8484 63812 10446
rect 63980 9938 64036 10556
rect 63980 9886 63982 9938
rect 64034 9886 64036 9938
rect 63980 9874 64036 9886
rect 64204 10498 64260 10510
rect 64204 10446 64206 10498
rect 64258 10446 64260 10498
rect 63756 8418 63812 8428
rect 63868 9268 63924 9278
rect 63868 8148 63924 9212
rect 64204 9268 64260 10446
rect 64204 9202 64260 9212
rect 64316 9602 64372 9614
rect 64316 9550 64318 9602
rect 64370 9550 64372 9602
rect 64204 8932 64260 8942
rect 64204 8838 64260 8876
rect 63868 8082 63924 8092
rect 64092 8818 64148 8830
rect 64092 8766 64094 8818
rect 64146 8766 64148 8818
rect 63868 7476 63924 7486
rect 63644 7422 63646 7474
rect 63698 7422 63700 7474
rect 63644 7410 63700 7422
rect 63756 7474 63924 7476
rect 63756 7422 63870 7474
rect 63922 7422 63924 7474
rect 63756 7420 63924 7422
rect 63532 7362 63588 7374
rect 63532 7310 63534 7362
rect 63586 7310 63588 7362
rect 63532 7028 63588 7310
rect 63532 6962 63588 6972
rect 63420 6626 63476 6636
rect 63420 6356 63476 6366
rect 63420 6018 63476 6300
rect 63420 5966 63422 6018
rect 63474 5966 63476 6018
rect 63420 5954 63476 5966
rect 63644 6020 63700 6030
rect 63644 5926 63700 5964
rect 63756 5794 63812 7420
rect 63868 7410 63924 7420
rect 64092 6356 64148 8766
rect 64316 6468 64372 9550
rect 64428 9044 64484 9054
rect 64428 8950 64484 8988
rect 64540 8820 64596 12236
rect 64764 12068 64820 12078
rect 65436 12068 65492 12078
rect 64764 12066 65044 12068
rect 64764 12014 64766 12066
rect 64818 12014 65044 12066
rect 64764 12012 65044 12014
rect 64764 12002 64820 12012
rect 64876 10724 64932 10734
rect 64764 10500 64820 10510
rect 64764 10164 64820 10444
rect 64764 10098 64820 10108
rect 64764 9940 64820 9950
rect 64876 9940 64932 10668
rect 64764 9938 64932 9940
rect 64764 9886 64766 9938
rect 64818 9886 64932 9938
rect 64764 9884 64932 9886
rect 64764 9874 64820 9884
rect 64428 8764 64596 8820
rect 64652 8820 64708 8830
rect 64428 8428 64484 8764
rect 64428 8372 64596 8428
rect 64316 6402 64372 6412
rect 64092 6290 64148 6300
rect 64316 6244 64372 6254
rect 64316 6018 64372 6188
rect 64316 5966 64318 6018
rect 64370 5966 64372 6018
rect 64316 5954 64372 5966
rect 63756 5742 63758 5794
rect 63810 5742 63812 5794
rect 63756 5730 63812 5742
rect 64428 5796 64484 5806
rect 64092 5010 64148 5022
rect 64092 4958 64094 5010
rect 64146 4958 64148 5010
rect 63644 4898 63700 4910
rect 63644 4846 63646 4898
rect 63698 4846 63700 4898
rect 63532 4450 63588 4462
rect 63532 4398 63534 4450
rect 63586 4398 63588 4450
rect 63532 3780 63588 4398
rect 63644 4116 63700 4846
rect 64092 4900 64148 4958
rect 64092 4834 64148 4844
rect 64316 5012 64372 5022
rect 64316 4562 64372 4956
rect 64428 5010 64484 5740
rect 64428 4958 64430 5010
rect 64482 4958 64484 5010
rect 64428 4946 64484 4958
rect 64316 4510 64318 4562
rect 64370 4510 64372 4562
rect 64316 4498 64372 4510
rect 64428 4788 64484 4798
rect 64428 4452 64484 4732
rect 64428 4358 64484 4396
rect 63644 4050 63700 4060
rect 64092 4338 64148 4350
rect 64092 4286 64094 4338
rect 64146 4286 64148 4338
rect 64092 4228 64148 4286
rect 64540 4228 64596 8372
rect 64652 7364 64708 8764
rect 64652 7362 64820 7364
rect 64652 7310 64654 7362
rect 64706 7310 64820 7362
rect 64652 7308 64820 7310
rect 64652 7298 64708 7308
rect 64652 6018 64708 6030
rect 64652 5966 64654 6018
rect 64706 5966 64708 6018
rect 64652 4452 64708 5966
rect 64652 4386 64708 4396
rect 64764 4228 64820 7308
rect 64876 6692 64932 9884
rect 64876 6626 64932 6636
rect 64988 5010 65044 12012
rect 65212 9604 65268 9614
rect 65100 6802 65156 6814
rect 65100 6750 65102 6802
rect 65154 6750 65156 6802
rect 65100 6020 65156 6750
rect 65212 6244 65268 9548
rect 65436 9604 65492 12012
rect 65548 10834 65604 24108
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 67004 19348 67060 19358
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65660 12066 65716 12078
rect 65660 12014 65662 12066
rect 65714 12014 65716 12066
rect 65660 11060 65716 12014
rect 66108 12068 66164 12078
rect 66108 11974 66164 12012
rect 66892 12068 66948 12078
rect 66892 11974 66948 12012
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 66556 11394 66612 11406
rect 66556 11342 66558 11394
rect 66610 11342 66612 11394
rect 65884 11284 65940 11294
rect 65884 11282 66500 11284
rect 65884 11230 65886 11282
rect 65938 11230 66500 11282
rect 65884 11228 66500 11230
rect 65884 11218 65940 11228
rect 65660 10994 65716 11004
rect 66332 11060 66388 11070
rect 65548 10782 65550 10834
rect 65602 10782 65604 10834
rect 65548 10500 65604 10782
rect 65548 10434 65604 10444
rect 65996 10724 66052 10734
rect 65996 10498 66052 10668
rect 65996 10446 65998 10498
rect 66050 10446 66052 10498
rect 65996 10434 66052 10446
rect 65916 10220 66180 10230
rect 65436 9510 65492 9548
rect 65548 10164 65604 10174
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 65436 9268 65492 9278
rect 65436 9174 65492 9212
rect 65212 6178 65268 6188
rect 65324 9156 65380 9166
rect 65100 5460 65156 5964
rect 65100 5394 65156 5404
rect 64988 4958 64990 5010
rect 65042 4958 65044 5010
rect 64092 4172 64596 4228
rect 64652 4172 64820 4228
rect 64876 4228 64932 4238
rect 63532 3714 63588 3724
rect 63532 3556 63588 3566
rect 63308 3554 63588 3556
rect 63308 3502 63534 3554
rect 63586 3502 63588 3554
rect 63308 3500 63588 3502
rect 63532 3490 63588 3500
rect 64092 980 64148 4172
rect 64316 3780 64372 3790
rect 64092 914 64148 924
rect 64204 3778 64372 3780
rect 64204 3726 64318 3778
rect 64370 3726 64372 3778
rect 64204 3724 64372 3726
rect 64204 800 64260 3724
rect 64316 3714 64372 3724
rect 64652 1092 64708 4172
rect 64764 4004 64820 4014
rect 64764 3668 64820 3948
rect 64764 3536 64820 3612
rect 64876 2100 64932 4172
rect 64988 3778 65044 4958
rect 65324 5010 65380 9100
rect 65548 6132 65604 10108
rect 65772 9940 65828 9950
rect 65772 9266 65828 9884
rect 65772 9214 65774 9266
rect 65826 9214 65828 9266
rect 65772 9202 65828 9214
rect 66220 9268 66276 9278
rect 66220 9174 66276 9212
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 66332 8428 66388 11004
rect 66444 9716 66500 11228
rect 66556 11172 66612 11342
rect 66556 9940 66612 11116
rect 66556 9874 66612 9884
rect 66444 9660 66836 9716
rect 66780 8930 66836 9660
rect 66892 9268 66948 9278
rect 66892 9174 66948 9212
rect 66780 8878 66782 8930
rect 66834 8878 66836 8930
rect 66780 8866 66836 8878
rect 67004 8428 67060 19292
rect 67340 12738 67396 12750
rect 67340 12686 67342 12738
rect 67394 12686 67396 12738
rect 67116 11172 67172 11182
rect 67116 11078 67172 11116
rect 67340 10724 67396 12686
rect 67452 12066 67508 12078
rect 67452 12014 67454 12066
rect 67506 12014 67508 12066
rect 67452 11060 67508 12014
rect 67452 10994 67508 11004
rect 67788 11508 67844 11518
rect 67900 11508 67956 27356
rect 68796 25396 68852 25406
rect 68236 19796 68292 19806
rect 68236 13074 68292 19740
rect 68796 13636 68852 25340
rect 69916 22708 69972 116172
rect 71372 116228 71428 116398
rect 69916 22642 69972 22652
rect 70140 28644 70196 28654
rect 69692 22148 69748 22158
rect 68796 13570 68852 13580
rect 69132 13636 69188 13646
rect 69132 13542 69188 13580
rect 69580 13636 69636 13646
rect 69580 13542 69636 13580
rect 68236 13022 68238 13074
rect 68290 13022 68292 13074
rect 68124 12066 68180 12078
rect 68124 12014 68126 12066
rect 68178 12014 68180 12066
rect 68124 11954 68180 12014
rect 68124 11902 68126 11954
rect 68178 11902 68180 11954
rect 68124 11890 68180 11902
rect 67788 11506 67956 11508
rect 67788 11454 67790 11506
rect 67842 11454 67956 11506
rect 67788 11452 67956 11454
rect 66332 8372 66612 8428
rect 66444 8148 66500 8158
rect 66444 7476 66500 8092
rect 66444 7410 66500 7420
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 65548 6000 65604 6076
rect 65660 6692 65716 6702
rect 65884 6692 65940 6702
rect 65716 6690 65940 6692
rect 65716 6638 65886 6690
rect 65938 6638 65940 6690
rect 65716 6636 65940 6638
rect 65436 5796 65492 5806
rect 65436 5702 65492 5740
rect 65324 4958 65326 5010
rect 65378 4958 65380 5010
rect 65324 4946 65380 4958
rect 65548 5460 65604 5470
rect 64988 3726 64990 3778
rect 65042 3726 65044 3778
rect 64988 3714 65044 3726
rect 65212 4676 65268 4686
rect 65212 3554 65268 4620
rect 65548 4338 65604 5404
rect 65660 5236 65716 6636
rect 65884 6626 65940 6636
rect 66108 6692 66164 6702
rect 65660 5170 65716 5180
rect 65772 6468 65828 6478
rect 65772 4900 65828 6412
rect 66108 6244 66164 6636
rect 66332 6690 66388 6702
rect 66332 6638 66334 6690
rect 66386 6638 66388 6690
rect 66332 6244 66388 6638
rect 66556 6690 66612 8372
rect 66892 8372 67060 8428
rect 67116 8818 67172 8830
rect 67116 8766 67118 8818
rect 67170 8766 67172 8818
rect 66892 7700 66948 8372
rect 66556 6638 66558 6690
rect 66610 6638 66612 6690
rect 66556 6468 66612 6638
rect 66556 6402 66612 6412
rect 66668 7644 66948 7700
rect 66556 6244 66612 6254
rect 66332 6188 66500 6244
rect 66108 6018 66164 6188
rect 66108 5966 66110 6018
rect 66162 5966 66164 6018
rect 66108 5954 66164 5966
rect 66332 6020 66388 6030
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 66332 5348 66388 5964
rect 66332 5122 66388 5292
rect 66332 5070 66334 5122
rect 66386 5070 66388 5122
rect 66332 5058 66388 5070
rect 65772 4834 65828 4844
rect 66444 4676 66500 6188
rect 66556 6130 66612 6188
rect 66556 6078 66558 6130
rect 66610 6078 66612 6130
rect 66556 6066 66612 6078
rect 66444 4610 66500 4620
rect 66668 5684 66724 7644
rect 66892 7476 66948 7486
rect 66892 7382 66948 7420
rect 66668 4676 66724 5628
rect 66780 6580 66836 6590
rect 66780 5906 66836 6524
rect 67004 6468 67060 6478
rect 67004 6374 67060 6412
rect 66780 5854 66782 5906
rect 66834 5854 66836 5906
rect 66780 5796 66836 5854
rect 66780 5122 66836 5740
rect 66780 5070 66782 5122
rect 66834 5070 66836 5122
rect 66780 5058 66836 5070
rect 67116 5124 67172 8766
rect 67340 8258 67396 10668
rect 67340 8206 67342 8258
rect 67394 8206 67396 8258
rect 67340 8194 67396 8206
rect 67564 10500 67620 10510
rect 67452 6356 67508 6366
rect 67228 6132 67284 6142
rect 67228 6018 67284 6076
rect 67228 5966 67230 6018
rect 67282 5966 67284 6018
rect 67228 5954 67284 5966
rect 67452 5906 67508 6300
rect 67564 6132 67620 10444
rect 67788 10276 67844 11452
rect 68124 11172 68180 11182
rect 68124 11078 68180 11116
rect 68124 10500 68180 10510
rect 67788 10210 67844 10220
rect 67900 10498 68180 10500
rect 67900 10446 68126 10498
rect 68178 10446 68180 10498
rect 67900 10444 68180 10446
rect 67676 9714 67732 9726
rect 67676 9662 67678 9714
rect 67730 9662 67732 9714
rect 67676 8932 67732 9662
rect 67788 9268 67844 9278
rect 67788 9174 67844 9212
rect 67900 9266 67956 10444
rect 68124 10434 68180 10444
rect 67900 9214 67902 9266
rect 67954 9214 67956 9266
rect 67900 9202 67956 9214
rect 68124 10276 68180 10286
rect 67676 8866 67732 8876
rect 68012 8818 68068 8830
rect 68012 8766 68014 8818
rect 68066 8766 68068 8818
rect 67676 8036 67732 8046
rect 67676 8034 67844 8036
rect 67676 7982 67678 8034
rect 67730 7982 67844 8034
rect 67676 7980 67844 7982
rect 67676 7970 67732 7980
rect 67788 6692 67844 7980
rect 68012 7140 68068 8766
rect 68124 8428 68180 10220
rect 68236 8708 68292 13022
rect 69692 13074 69748 22092
rect 69692 13022 69694 13074
rect 69746 13022 69748 13074
rect 68460 12852 68516 12862
rect 68460 12404 68516 12796
rect 68684 12740 68740 12750
rect 68348 9828 68404 9838
rect 68348 9734 68404 9772
rect 68236 8642 68292 8652
rect 68124 8372 68292 8428
rect 68236 8370 68292 8372
rect 68236 8318 68238 8370
rect 68290 8318 68292 8370
rect 68236 8306 68292 8318
rect 68012 7074 68068 7084
rect 68124 6692 68180 6702
rect 67788 6636 68068 6692
rect 67676 6580 67732 6590
rect 67676 6486 67732 6524
rect 67900 6466 67956 6478
rect 67900 6414 67902 6466
rect 67954 6414 67956 6466
rect 67676 6132 67732 6142
rect 67564 6130 67732 6132
rect 67564 6078 67678 6130
rect 67730 6078 67732 6130
rect 67564 6076 67732 6078
rect 67676 6066 67732 6076
rect 67788 6132 67844 6142
rect 67788 6038 67844 6076
rect 67900 6020 67956 6414
rect 67900 5954 67956 5964
rect 67452 5854 67454 5906
rect 67506 5854 67508 5906
rect 67452 5684 67508 5854
rect 67564 5908 67620 5918
rect 67564 5814 67620 5852
rect 67508 5628 67620 5684
rect 67452 5618 67508 5628
rect 67116 5068 67508 5124
rect 66892 5012 66948 5022
rect 66892 5010 67396 5012
rect 66892 4958 66894 5010
rect 66946 4958 67396 5010
rect 66892 4956 67396 4958
rect 66892 4946 66948 4956
rect 66668 4610 66724 4620
rect 65548 4286 65550 4338
rect 65602 4286 65604 4338
rect 65548 4274 65604 4286
rect 67340 4338 67396 4956
rect 67452 4900 67508 5068
rect 67452 4834 67508 4844
rect 67564 4452 67620 5628
rect 67676 5124 67732 5134
rect 67676 5030 67732 5068
rect 67788 4900 67844 4910
rect 67788 4562 67844 4844
rect 68012 4900 68068 6636
rect 68460 6692 68516 12348
rect 68572 12738 68740 12740
rect 68572 12686 68686 12738
rect 68738 12686 68740 12738
rect 68572 12684 68740 12686
rect 68572 11954 68628 12684
rect 68684 12674 68740 12684
rect 68684 12068 68740 12078
rect 69132 12068 69188 12078
rect 69580 12068 69636 12078
rect 68684 12066 69636 12068
rect 68684 12014 68686 12066
rect 68738 12014 69134 12066
rect 69186 12014 69582 12066
rect 69634 12014 69636 12066
rect 68684 12012 69636 12014
rect 68684 12002 68740 12012
rect 69132 12002 69188 12012
rect 68572 11902 68574 11954
rect 68626 11902 68628 11954
rect 68572 11396 68628 11902
rect 68572 11330 68628 11340
rect 69132 11732 69188 11742
rect 68572 11172 68628 11182
rect 68572 11078 68628 11116
rect 68684 11060 68740 11070
rect 68572 10948 68628 10958
rect 68572 9492 68628 10892
rect 68572 9426 68628 9436
rect 68684 9268 68740 11004
rect 68796 10610 68852 10622
rect 68796 10558 68798 10610
rect 68850 10558 68852 10610
rect 68796 9828 68852 10558
rect 68852 9772 69076 9828
rect 68796 9762 68852 9772
rect 68684 9136 68740 9212
rect 68796 9492 68852 9502
rect 68796 9044 68852 9436
rect 68684 8988 68852 9044
rect 69020 9044 69076 9772
rect 68572 8932 68628 8942
rect 68572 8838 68628 8876
rect 68572 8372 68628 8382
rect 68684 8372 68740 8988
rect 68908 8818 68964 8830
rect 68908 8766 68910 8818
rect 68962 8766 68964 8818
rect 68572 8370 68740 8372
rect 68572 8318 68574 8370
rect 68626 8318 68740 8370
rect 68572 8316 68740 8318
rect 68796 8708 68852 8718
rect 68572 8306 68628 8316
rect 68572 6692 68628 6702
rect 68460 6690 68628 6692
rect 68460 6638 68574 6690
rect 68626 6638 68628 6690
rect 68460 6636 68628 6638
rect 68124 6578 68180 6636
rect 68572 6626 68628 6636
rect 68124 6526 68126 6578
rect 68178 6526 68180 6578
rect 68124 6514 68180 6526
rect 68236 6466 68292 6478
rect 68236 6414 68238 6466
rect 68290 6414 68292 6466
rect 68236 5236 68292 6414
rect 68796 6132 68852 8652
rect 68908 7252 68964 8766
rect 69020 7586 69076 8988
rect 69020 7534 69022 7586
rect 69074 7534 69076 7586
rect 69020 7522 69076 7534
rect 69132 7252 69188 11676
rect 69244 11172 69300 11182
rect 69244 11078 69300 11116
rect 68908 7186 68964 7196
rect 69020 7196 69188 7252
rect 69244 10612 69300 10622
rect 68796 6066 68852 6076
rect 68460 5906 68516 5918
rect 68460 5854 68462 5906
rect 68514 5854 68516 5906
rect 68460 5346 68516 5854
rect 68796 5906 68852 5918
rect 68796 5854 68798 5906
rect 68850 5854 68852 5906
rect 68796 5684 68852 5854
rect 69020 5908 69076 7196
rect 69132 5908 69188 5918
rect 69020 5906 69188 5908
rect 69020 5854 69134 5906
rect 69186 5854 69188 5906
rect 69020 5852 69188 5854
rect 69132 5842 69188 5852
rect 68796 5618 68852 5628
rect 68908 5684 68964 5694
rect 69244 5684 69300 10556
rect 69356 9826 69412 12012
rect 69580 12002 69636 12012
rect 69692 11732 69748 13022
rect 70028 13634 70084 13646
rect 70028 13582 70030 13634
rect 70082 13582 70084 13634
rect 69692 11666 69748 11676
rect 69804 12068 69860 12078
rect 69692 11396 69748 11406
rect 69692 11302 69748 11340
rect 69692 10500 69748 10510
rect 69804 10500 69860 12012
rect 70028 12068 70084 13582
rect 70140 13076 70196 28588
rect 71372 27412 71428 116172
rect 72268 116228 72324 116238
rect 72268 116134 72324 116172
rect 72604 115556 72660 115566
rect 72604 115462 72660 115500
rect 71372 27346 71428 27356
rect 72156 25284 72212 25294
rect 70140 12944 70196 13020
rect 70252 24052 70308 24062
rect 70252 12404 70308 23996
rect 71260 20580 71316 20590
rect 70588 13636 70644 13646
rect 70588 13634 70756 13636
rect 70588 13582 70590 13634
rect 70642 13582 70756 13634
rect 70588 13580 70756 13582
rect 70588 13570 70644 13580
rect 70252 12272 70308 12348
rect 70028 12002 70084 12012
rect 70588 12068 70644 12078
rect 70588 11974 70644 12012
rect 70700 11620 70756 13580
rect 71036 13634 71092 13646
rect 71036 13582 71038 13634
rect 71090 13582 71092 13634
rect 71036 12964 71092 13582
rect 71036 12898 71092 12908
rect 71260 13074 71316 20524
rect 71260 13022 71262 13074
rect 71314 13022 71316 13074
rect 70812 12740 70868 12750
rect 70812 12738 71204 12740
rect 70812 12686 70814 12738
rect 70866 12686 71204 12738
rect 70812 12684 71204 12686
rect 70812 12674 70868 12684
rect 70924 12516 70980 12526
rect 70700 11564 70868 11620
rect 70140 11508 70196 11518
rect 70812 11508 70868 11564
rect 70196 11452 70308 11508
rect 70140 11414 70196 11452
rect 69692 10498 69860 10500
rect 69692 10446 69694 10498
rect 69746 10446 69860 10498
rect 69692 10444 69860 10446
rect 69692 10434 69748 10444
rect 69356 9774 69358 9826
rect 69410 9774 69412 9826
rect 69356 8258 69412 9774
rect 69692 8932 69748 8942
rect 69692 8838 69748 8876
rect 69804 8428 69860 10444
rect 69356 8206 69358 8258
rect 69410 8206 69412 8258
rect 69356 7476 69412 8206
rect 69468 8372 69860 8428
rect 70028 11396 70084 11406
rect 70028 8596 70084 11340
rect 69468 8148 69524 8372
rect 69468 8082 69524 8092
rect 69356 6690 69412 7420
rect 69804 7364 69860 7374
rect 69692 7252 69748 7262
rect 69356 6638 69358 6690
rect 69410 6638 69412 6690
rect 69356 6626 69412 6638
rect 69468 7140 69524 7150
rect 69468 6130 69524 7084
rect 69468 6078 69470 6130
rect 69522 6078 69524 6130
rect 69468 6066 69524 6078
rect 69356 6020 69412 6030
rect 69356 5926 69412 5964
rect 68908 5682 69300 5684
rect 68908 5630 68910 5682
rect 68962 5630 69300 5682
rect 68908 5628 69300 5630
rect 68908 5618 68964 5628
rect 68460 5294 68462 5346
rect 68514 5294 68516 5346
rect 68460 5282 68516 5294
rect 68236 5104 68292 5180
rect 69580 5236 69636 5246
rect 68012 4834 68068 4844
rect 69356 5010 69412 5022
rect 69356 4958 69358 5010
rect 69410 4958 69412 5010
rect 69356 4788 69412 4958
rect 69580 5010 69636 5180
rect 69580 4958 69582 5010
rect 69634 4958 69636 5010
rect 69580 4946 69636 4958
rect 69692 4898 69748 7196
rect 69804 5346 69860 7308
rect 70028 6468 70084 8540
rect 70028 5906 70084 6412
rect 70028 5854 70030 5906
rect 70082 5854 70084 5906
rect 70028 5842 70084 5854
rect 70140 10948 70196 10958
rect 69804 5294 69806 5346
rect 69858 5294 69860 5346
rect 69804 5282 69860 5294
rect 70028 5236 70084 5246
rect 70140 5236 70196 10892
rect 70252 10836 70308 11452
rect 70700 11396 70756 11406
rect 70700 11302 70756 11340
rect 70812 11282 70868 11452
rect 70812 11230 70814 11282
rect 70866 11230 70868 11282
rect 70812 11218 70868 11230
rect 70252 8428 70308 10780
rect 70812 8596 70868 8606
rect 70252 8372 70532 8428
rect 70252 5906 70308 8372
rect 70252 5854 70254 5906
rect 70306 5854 70308 5906
rect 70252 5842 70308 5854
rect 70028 5234 70196 5236
rect 70028 5182 70030 5234
rect 70082 5182 70196 5234
rect 70028 5180 70196 5182
rect 70028 5170 70084 5180
rect 70252 5124 70308 5134
rect 70252 5030 70308 5068
rect 70476 5012 70532 8372
rect 70476 4946 70532 4956
rect 70588 6244 70644 6254
rect 69692 4846 69694 4898
rect 69746 4846 69748 4898
rect 69692 4834 69748 4846
rect 70364 4900 70420 4910
rect 69356 4722 69412 4732
rect 67788 4510 67790 4562
rect 67842 4510 67844 4562
rect 67788 4498 67844 4510
rect 68124 4676 68180 4686
rect 67676 4452 67732 4462
rect 67564 4450 67732 4452
rect 67564 4398 67678 4450
rect 67730 4398 67732 4450
rect 67564 4396 67732 4398
rect 67676 4386 67732 4396
rect 67900 4452 67956 4462
rect 67340 4286 67342 4338
rect 67394 4286 67396 4338
rect 67340 4274 67396 4286
rect 67900 4338 67956 4396
rect 67900 4286 67902 4338
rect 67954 4286 67956 4338
rect 67900 4274 67956 4286
rect 68124 4338 68180 4620
rect 68908 4676 68964 4686
rect 68908 4562 68964 4620
rect 68908 4510 68910 4562
rect 68962 4510 68964 4562
rect 68908 4498 68964 4510
rect 68348 4452 68404 4462
rect 68348 4358 68404 4396
rect 68124 4286 68126 4338
rect 68178 4286 68180 4338
rect 68124 4274 68180 4286
rect 69356 4340 69412 4350
rect 69356 4246 69412 4284
rect 66108 4228 66164 4238
rect 66108 4134 66164 4172
rect 69244 4228 69300 4238
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 66108 3780 66164 3790
rect 65212 3502 65214 3554
rect 65266 3502 65268 3554
rect 65212 3490 65268 3502
rect 65548 3556 65604 3566
rect 65548 3330 65604 3500
rect 66108 3554 66164 3724
rect 66108 3502 66110 3554
rect 66162 3502 66164 3554
rect 66108 3490 66164 3502
rect 68460 3556 68516 3566
rect 68460 3462 68516 3500
rect 65548 3278 65550 3330
rect 65602 3278 65604 3330
rect 65548 3266 65604 3278
rect 65884 3444 65940 3454
rect 64652 1026 64708 1036
rect 64764 2044 64932 2100
rect 64764 800 64820 2044
rect 65884 800 65940 3388
rect 67004 3444 67060 3454
rect 67004 3350 67060 3388
rect 67564 3444 67620 3454
rect 67564 800 67620 3388
rect 69244 800 69300 4172
rect 70028 4228 70084 4238
rect 70028 4134 70084 4172
rect 70364 3554 70420 4844
rect 70588 4788 70644 6188
rect 70588 4722 70644 4732
rect 70700 5908 70756 5918
rect 70364 3502 70366 3554
rect 70418 3502 70420 3554
rect 70364 3490 70420 3502
rect 69356 3444 69412 3454
rect 69356 3350 69412 3388
rect 70700 1204 70756 5852
rect 70812 5010 70868 8540
rect 70924 6468 70980 12460
rect 71036 12068 71092 12078
rect 71036 11844 71092 12012
rect 71036 11778 71092 11788
rect 71036 11170 71092 11182
rect 71036 11118 71038 11170
rect 71090 11118 71092 11170
rect 71036 7364 71092 11118
rect 71148 10612 71204 12684
rect 71260 10948 71316 13022
rect 71260 10882 71316 10892
rect 71372 13636 71428 13646
rect 71148 10556 71316 10612
rect 71036 7298 71092 7308
rect 71148 10388 71204 10398
rect 70924 6402 70980 6412
rect 70812 4958 70814 5010
rect 70866 4958 70868 5010
rect 70812 4900 70868 4958
rect 70812 4834 70868 4844
rect 70924 5794 70980 5806
rect 70924 5742 70926 5794
rect 70978 5742 70980 5794
rect 70924 4452 70980 5742
rect 71036 5012 71092 5022
rect 71036 4918 71092 4956
rect 70924 4386 70980 4396
rect 71148 4338 71204 10332
rect 71260 10052 71316 10556
rect 71260 9986 71316 9996
rect 71260 8148 71316 8158
rect 71260 7476 71316 8092
rect 71260 7028 71316 7420
rect 71260 5012 71316 6972
rect 71372 5684 71428 13580
rect 72156 13076 72212 25228
rect 72940 15316 72996 15326
rect 72716 13636 72772 13646
rect 72716 13542 72772 13580
rect 72268 13076 72324 13086
rect 72156 13074 72324 13076
rect 72156 13022 72270 13074
rect 72322 13022 72324 13074
rect 72156 13020 72324 13022
rect 71484 12964 71540 12974
rect 71484 10836 71540 12908
rect 71708 12738 71764 12750
rect 71708 12686 71710 12738
rect 71762 12686 71764 12738
rect 71596 11732 71652 11742
rect 71596 11172 71652 11676
rect 71708 11396 71764 12686
rect 72156 12516 72212 13020
rect 72268 13010 72324 13020
rect 72156 12450 72212 12460
rect 72716 12738 72772 12750
rect 72716 12686 72718 12738
rect 72770 12686 72772 12738
rect 72268 12404 72324 12414
rect 71932 12066 71988 12078
rect 71932 12014 71934 12066
rect 71986 12014 71988 12066
rect 71932 11732 71988 12014
rect 71932 11666 71988 11676
rect 71708 11330 71764 11340
rect 71820 11284 71876 11294
rect 71820 11282 72212 11284
rect 71820 11230 71822 11282
rect 71874 11230 72212 11282
rect 71820 11228 72212 11230
rect 71820 11218 71876 11228
rect 71596 11078 71652 11116
rect 71708 11170 71764 11182
rect 71708 11118 71710 11170
rect 71762 11118 71764 11170
rect 71484 10770 71540 10780
rect 71708 9156 71764 11118
rect 71820 10498 71876 10510
rect 71820 10446 71822 10498
rect 71874 10446 71876 10498
rect 71820 10164 71876 10446
rect 71820 10098 71876 10108
rect 71932 10052 71988 10062
rect 71820 9156 71876 9166
rect 71708 9154 71876 9156
rect 71708 9102 71822 9154
rect 71874 9102 71876 9154
rect 71708 9100 71876 9102
rect 71820 9090 71876 9100
rect 71596 7476 71652 7486
rect 71596 7382 71652 7420
rect 71708 7364 71764 7374
rect 71708 7270 71764 7308
rect 71932 6244 71988 9996
rect 71932 6178 71988 6188
rect 72044 6468 72100 6478
rect 71932 5906 71988 5918
rect 71932 5854 71934 5906
rect 71986 5854 71988 5906
rect 71372 5618 71428 5628
rect 71820 5794 71876 5806
rect 71820 5742 71822 5794
rect 71874 5742 71876 5794
rect 71820 5460 71876 5742
rect 71372 5404 71876 5460
rect 71372 5346 71428 5404
rect 71372 5294 71374 5346
rect 71426 5294 71428 5346
rect 71372 5282 71428 5294
rect 71932 5348 71988 5854
rect 71932 5282 71988 5292
rect 71260 4918 71316 4956
rect 71708 5236 71764 5246
rect 71372 4564 71428 4574
rect 71372 4470 71428 4508
rect 71148 4286 71150 4338
rect 71202 4286 71204 4338
rect 71148 4274 71204 4286
rect 71708 4338 71764 5180
rect 71820 4452 71876 4462
rect 71820 4358 71876 4396
rect 71708 4286 71710 4338
rect 71762 4286 71764 4338
rect 71708 4274 71764 4286
rect 72044 4226 72100 6412
rect 72156 4562 72212 11228
rect 72268 8932 72324 12348
rect 72380 12066 72436 12078
rect 72380 12014 72382 12066
rect 72434 12014 72436 12066
rect 72380 11396 72436 12014
rect 72604 11396 72660 11406
rect 72380 11394 72660 11396
rect 72380 11342 72606 11394
rect 72658 11342 72660 11394
rect 72380 11340 72660 11342
rect 72492 10612 72548 10622
rect 72604 10612 72660 11340
rect 72492 10610 72660 10612
rect 72492 10558 72494 10610
rect 72546 10558 72660 10610
rect 72492 10556 72660 10558
rect 72492 9044 72548 10556
rect 72716 9380 72772 12686
rect 72716 9314 72772 9324
rect 72492 8950 72548 8988
rect 72268 6132 72324 8876
rect 72268 5122 72324 6076
rect 72380 7250 72436 7262
rect 72380 7198 72382 7250
rect 72434 7198 72436 7250
rect 72380 6020 72436 7198
rect 72380 5954 72436 5964
rect 72268 5070 72270 5122
rect 72322 5070 72324 5122
rect 72268 5058 72324 5070
rect 72604 5906 72660 5918
rect 72604 5854 72606 5906
rect 72658 5854 72660 5906
rect 72492 5010 72548 5022
rect 72492 4958 72494 5010
rect 72546 4958 72548 5010
rect 72492 4900 72548 4958
rect 72492 4834 72548 4844
rect 72156 4510 72158 4562
rect 72210 4510 72212 4562
rect 72156 4498 72212 4510
rect 72604 4452 72660 5854
rect 72604 4386 72660 4396
rect 72380 4340 72436 4350
rect 72380 4246 72436 4284
rect 72940 4340 72996 15260
rect 73052 12068 73108 116508
rect 73500 116564 73556 119200
rect 73500 116498 73556 116508
rect 74396 116564 74452 116574
rect 74396 116470 74452 116508
rect 75068 116564 75124 119200
rect 77532 117010 77588 117022
rect 77532 116958 77534 117010
rect 77586 116958 77588 117010
rect 75068 116498 75124 116508
rect 76524 116564 76580 116574
rect 76524 116470 76580 116508
rect 73724 116450 73780 116462
rect 73724 116398 73726 116450
rect 73778 116398 73780 116450
rect 73724 115890 73780 116398
rect 77532 116450 77588 116958
rect 78204 116676 78260 119200
rect 78204 116610 78260 116620
rect 78652 117010 78708 117022
rect 78652 116958 78654 117010
rect 78706 116958 78708 117010
rect 77532 116398 77534 116450
rect 77586 116398 77588 116450
rect 77532 116386 77588 116398
rect 78204 116450 78260 116462
rect 78204 116398 78206 116450
rect 78258 116398 78260 116450
rect 73724 115838 73726 115890
rect 73778 115838 73780 115890
rect 73724 115826 73780 115838
rect 78204 115890 78260 116398
rect 78204 115838 78206 115890
rect 78258 115838 78260 115890
rect 78204 115826 78260 115838
rect 78652 115890 78708 116958
rect 78988 116676 79044 116686
rect 78988 116562 79044 116620
rect 78988 116510 78990 116562
rect 79042 116510 79044 116562
rect 78988 116498 79044 116510
rect 79772 116564 79828 119200
rect 79772 116498 79828 116508
rect 80668 116564 80724 116574
rect 80668 116470 80724 116508
rect 81228 116452 81284 116462
rect 81900 116452 81956 116462
rect 81116 116450 81956 116452
rect 81116 116398 81230 116450
rect 81282 116398 81902 116450
rect 81954 116398 81956 116450
rect 81116 116396 81956 116398
rect 78652 115838 78654 115890
rect 78706 115838 78708 115890
rect 73500 115666 73556 115678
rect 73500 115614 73502 115666
rect 73554 115614 73556 115666
rect 73500 115556 73556 115614
rect 77980 115666 78036 115678
rect 77980 115614 77982 115666
rect 78034 115614 78036 115666
rect 73500 115490 73556 115500
rect 77308 115556 77364 115566
rect 77308 115462 77364 115500
rect 77980 115556 78036 115614
rect 77980 115490 78036 115500
rect 74844 29428 74900 29438
rect 74732 22484 74788 22494
rect 73948 22260 74004 22270
rect 73948 13524 74004 22204
rect 73500 13468 73948 13524
rect 73500 13074 73556 13468
rect 73948 13458 74004 13468
rect 74060 14420 74116 14430
rect 73500 13022 73502 13074
rect 73554 13022 73556 13074
rect 73500 13010 73556 13022
rect 73052 12002 73108 12012
rect 73164 12738 73220 12750
rect 73164 12686 73166 12738
rect 73218 12686 73220 12738
rect 73164 5908 73220 12686
rect 73612 12292 73668 12302
rect 73668 12236 73892 12292
rect 73612 12198 73668 12236
rect 73388 11396 73444 11406
rect 73388 11394 73668 11396
rect 73388 11342 73390 11394
rect 73442 11342 73668 11394
rect 73388 11340 73668 11342
rect 73388 11330 73444 11340
rect 73276 11172 73332 11182
rect 73276 10388 73332 11116
rect 73500 11172 73556 11182
rect 73388 10612 73444 10622
rect 73388 10518 73444 10556
rect 73276 10332 73444 10388
rect 73164 5842 73220 5852
rect 73276 9380 73332 9390
rect 73276 4340 73332 9324
rect 73388 7698 73444 10332
rect 73500 8370 73556 11116
rect 73612 8930 73668 11340
rect 73836 10836 73892 12236
rect 73724 10724 73780 10734
rect 73836 10724 73892 10780
rect 73948 10724 74004 10734
rect 73836 10722 74004 10724
rect 73836 10670 73950 10722
rect 74002 10670 74004 10722
rect 73836 10668 74004 10670
rect 73724 9716 73780 10668
rect 73948 10658 74004 10668
rect 73836 10500 73892 10510
rect 73836 9938 73892 10444
rect 73836 9886 73838 9938
rect 73890 9886 73892 9938
rect 73836 9874 73892 9886
rect 73724 9660 73892 9716
rect 73724 9268 73780 9278
rect 73724 9174 73780 9212
rect 73836 9044 73892 9660
rect 73612 8878 73614 8930
rect 73666 8878 73668 8930
rect 73612 8866 73668 8878
rect 73724 8988 73892 9044
rect 74060 9044 74116 14364
rect 74172 12738 74228 12750
rect 74732 12740 74788 22428
rect 74844 13076 74900 29372
rect 74956 22372 75012 22382
rect 74956 13636 75012 22316
rect 76076 21028 76132 21038
rect 74956 13634 75124 13636
rect 74956 13582 74958 13634
rect 75010 13582 75124 13634
rect 74956 13580 75124 13582
rect 74956 13570 75012 13580
rect 74844 13010 74900 13020
rect 74172 12686 74174 12738
rect 74226 12686 74228 12738
rect 74172 12404 74228 12686
rect 74172 12338 74228 12348
rect 74396 12738 74788 12740
rect 74396 12686 74734 12738
rect 74786 12686 74788 12738
rect 74396 12684 74788 12686
rect 74172 12066 74228 12078
rect 74172 12014 74174 12066
rect 74226 12014 74228 12066
rect 74172 11508 74228 12014
rect 74172 10836 74228 11452
rect 74284 10836 74340 10846
rect 74172 10834 74340 10836
rect 74172 10782 74286 10834
rect 74338 10782 74340 10834
rect 74172 10780 74340 10782
rect 74172 10724 74228 10780
rect 74284 10770 74340 10780
rect 74172 10658 74228 10668
rect 73500 8318 73502 8370
rect 73554 8318 73556 8370
rect 73500 8306 73556 8318
rect 73388 7646 73390 7698
rect 73442 7646 73444 7698
rect 73388 7634 73444 7646
rect 73724 7586 73780 8988
rect 74060 8978 74116 8988
rect 73948 8820 74004 8830
rect 73948 8818 74228 8820
rect 73948 8766 73950 8818
rect 74002 8766 74228 8818
rect 73948 8764 74228 8766
rect 73948 8754 74004 8764
rect 73724 7534 73726 7586
rect 73778 7534 73780 7586
rect 73724 7522 73780 7534
rect 73836 8484 73892 8494
rect 73836 6802 73892 8428
rect 73836 6750 73838 6802
rect 73890 6750 73892 6802
rect 73836 6738 73892 6750
rect 74060 6020 74116 6030
rect 74060 5926 74116 5964
rect 73388 5908 73444 5918
rect 73388 5814 73444 5852
rect 73612 5906 73668 5918
rect 73948 5908 74004 5918
rect 73612 5854 73614 5906
rect 73666 5854 73668 5906
rect 73612 5348 73668 5854
rect 73388 5292 73668 5348
rect 73724 5852 73948 5908
rect 73388 4788 73444 5292
rect 73500 5124 73556 5134
rect 73500 5010 73556 5068
rect 73500 4958 73502 5010
rect 73554 4958 73556 5010
rect 73500 4946 73556 4958
rect 73612 5122 73668 5134
rect 73612 5070 73614 5122
rect 73666 5070 73668 5122
rect 73612 5012 73668 5070
rect 73612 4946 73668 4956
rect 73388 4732 73668 4788
rect 73612 4564 73668 4732
rect 73388 4340 73444 4350
rect 73276 4338 73444 4340
rect 73276 4286 73390 4338
rect 73442 4286 73444 4338
rect 73276 4284 73444 4286
rect 72940 4274 72996 4284
rect 73388 4274 73444 4284
rect 73612 4338 73668 4508
rect 73612 4286 73614 4338
rect 73666 4286 73668 4338
rect 72044 4174 72046 4226
rect 72098 4174 72100 4226
rect 72044 4162 72100 4174
rect 71036 3668 71092 3678
rect 72716 3668 72772 3678
rect 70700 1138 70756 1148
rect 70924 3666 71092 3668
rect 70924 3614 71038 3666
rect 71090 3614 71092 3666
rect 70924 3612 71092 3614
rect 70924 800 70980 3612
rect 71036 3602 71092 3612
rect 72604 3666 72772 3668
rect 72604 3614 72718 3666
rect 72770 3614 72772 3666
rect 72604 3612 72772 3614
rect 72604 800 72660 3612
rect 72716 3602 72772 3612
rect 73612 3668 73668 4286
rect 73724 4338 73780 5852
rect 73948 5814 74004 5852
rect 73724 4286 73726 4338
rect 73778 4286 73780 4338
rect 73724 4274 73780 4286
rect 73836 5124 73892 5134
rect 73612 3602 73668 3612
rect 73724 3556 73780 3566
rect 73836 3556 73892 5068
rect 74172 4562 74228 8764
rect 74172 4510 74174 4562
rect 74226 4510 74228 4562
rect 74172 4498 74228 4510
rect 74284 7586 74340 7598
rect 74284 7534 74286 7586
rect 74338 7534 74340 7586
rect 74060 4452 74116 4462
rect 74060 4358 74116 4396
rect 73724 3554 73892 3556
rect 73724 3502 73726 3554
rect 73778 3502 73892 3554
rect 73724 3500 73892 3502
rect 74284 3554 74340 7534
rect 74396 5906 74452 12684
rect 74732 12674 74788 12684
rect 74956 12516 75012 12526
rect 74508 12066 74564 12078
rect 74508 12014 74510 12066
rect 74562 12014 74564 12066
rect 74508 11844 74564 12014
rect 74508 11778 74564 11788
rect 74956 12066 75012 12460
rect 74956 12014 74958 12066
rect 75010 12014 75012 12066
rect 74956 10948 75012 12014
rect 74508 10892 75012 10948
rect 74508 9268 74564 10892
rect 74956 10724 75012 10734
rect 74956 10630 75012 10668
rect 74844 10612 74900 10622
rect 74732 9716 74788 9726
rect 74620 9268 74676 9278
rect 74508 9266 74676 9268
rect 74508 9214 74622 9266
rect 74674 9214 74676 9266
rect 74508 9212 74676 9214
rect 74620 9202 74676 9212
rect 74508 9042 74564 9054
rect 74508 8990 74510 9042
rect 74562 8990 74564 9042
rect 74508 8260 74564 8990
rect 74620 9044 74676 9054
rect 74620 8818 74676 8988
rect 74620 8766 74622 8818
rect 74674 8766 74676 8818
rect 74620 8754 74676 8766
rect 74508 8194 74564 8204
rect 74508 7476 74564 7486
rect 74508 7382 74564 7420
rect 74732 6130 74788 9660
rect 74732 6078 74734 6130
rect 74786 6078 74788 6130
rect 74732 6066 74788 6078
rect 74396 5854 74398 5906
rect 74450 5854 74452 5906
rect 74396 5842 74452 5854
rect 74732 5796 74788 5806
rect 74396 4340 74452 4350
rect 74396 4246 74452 4284
rect 74284 3502 74286 3554
rect 74338 3502 74340 3554
rect 73724 3490 73780 3500
rect 74284 3490 74340 3502
rect 74620 4226 74676 4238
rect 74620 4174 74622 4226
rect 74674 4174 74676 4226
rect 74620 4116 74676 4174
rect 74396 3444 74452 3454
rect 74396 1764 74452 3388
rect 74620 2660 74676 4060
rect 74620 2594 74676 2604
rect 74732 2548 74788 5740
rect 74844 3892 74900 10556
rect 75068 10500 75124 13580
rect 75404 13634 75460 13646
rect 75852 13636 75908 13646
rect 75404 13582 75406 13634
rect 75458 13582 75460 13634
rect 75404 13524 75460 13582
rect 75404 13458 75460 13468
rect 75628 13634 75908 13636
rect 75628 13582 75854 13634
rect 75906 13582 75908 13634
rect 75628 13580 75908 13582
rect 75628 13524 75684 13580
rect 75852 13570 75908 13580
rect 75180 12740 75236 12750
rect 75180 12646 75236 12684
rect 75516 12066 75572 12078
rect 75516 12014 75518 12066
rect 75570 12014 75572 12066
rect 74956 10444 75124 10500
rect 75180 10610 75236 10622
rect 75180 10558 75182 10610
rect 75234 10558 75236 10610
rect 74956 4340 75012 10444
rect 75180 9940 75236 10558
rect 75068 9884 75236 9940
rect 75292 10164 75348 10174
rect 75292 9938 75348 10108
rect 75292 9886 75294 9938
rect 75346 9886 75348 9938
rect 75068 7476 75124 9884
rect 75292 9874 75348 9886
rect 75180 9716 75236 9726
rect 75180 9622 75236 9660
rect 75404 9602 75460 9614
rect 75404 9550 75406 9602
rect 75458 9550 75460 9602
rect 75292 9492 75348 9502
rect 75292 8372 75348 9436
rect 75404 9268 75460 9550
rect 75404 9202 75460 9212
rect 75404 9044 75460 9054
rect 75516 9044 75572 12014
rect 75460 8988 75572 9044
rect 75628 11170 75684 13468
rect 75740 13186 75796 13198
rect 75740 13134 75742 13186
rect 75794 13134 75796 13186
rect 75740 13074 75796 13134
rect 75740 13022 75742 13074
rect 75794 13022 75796 13074
rect 75740 13010 75796 13022
rect 75964 12852 76020 12862
rect 75852 12404 75908 12414
rect 75628 11118 75630 11170
rect 75682 11118 75684 11170
rect 75404 8484 75460 8988
rect 75404 8418 75460 8428
rect 75292 8260 75348 8316
rect 75516 8372 75572 8382
rect 75404 8260 75460 8270
rect 75292 8258 75460 8260
rect 75292 8206 75406 8258
rect 75458 8206 75460 8258
rect 75292 8204 75460 8206
rect 75404 8194 75460 8204
rect 75516 8146 75572 8316
rect 75516 8094 75518 8146
rect 75570 8094 75572 8146
rect 75516 7812 75572 8094
rect 75404 7700 75460 7710
rect 75404 7606 75460 7644
rect 75516 7588 75572 7756
rect 75516 7522 75572 7532
rect 75292 7476 75348 7486
rect 75068 7420 75292 7476
rect 75292 7382 75348 7420
rect 75292 7252 75348 7262
rect 75180 6468 75236 6478
rect 75068 6466 75236 6468
rect 75068 6414 75182 6466
rect 75234 6414 75236 6466
rect 75068 6412 75236 6414
rect 75068 5460 75124 6412
rect 75180 6402 75236 6412
rect 75068 5394 75124 5404
rect 75180 6018 75236 6030
rect 75180 5966 75182 6018
rect 75234 5966 75236 6018
rect 75180 5124 75236 5966
rect 75292 5684 75348 7196
rect 75404 7252 75460 7262
rect 75628 7252 75684 11118
rect 75740 12068 75796 12078
rect 75740 11396 75796 12012
rect 75740 10834 75796 11340
rect 75740 10782 75742 10834
rect 75794 10782 75796 10834
rect 75740 10770 75796 10782
rect 75852 8372 75908 12348
rect 75964 8932 76020 12796
rect 76076 12404 76132 20972
rect 77868 20804 77924 20814
rect 77644 15876 77700 15886
rect 77644 15148 77700 15820
rect 77532 15092 77700 15148
rect 77308 13860 77364 13870
rect 77084 13636 77140 13646
rect 76412 13186 76468 13198
rect 76412 13134 76414 13186
rect 76466 13134 76468 13186
rect 76076 12272 76132 12348
rect 76188 12738 76244 12750
rect 76188 12686 76190 12738
rect 76242 12686 76244 12738
rect 76188 12628 76244 12686
rect 76188 12180 76244 12572
rect 76188 12114 76244 12124
rect 76188 11170 76244 11182
rect 76188 11118 76190 11170
rect 76242 11118 76244 11170
rect 76188 11060 76244 11118
rect 76188 10724 76244 11004
rect 76188 10658 76244 10668
rect 76188 10500 76244 10510
rect 76188 10406 76244 10444
rect 76188 9938 76244 9950
rect 76188 9886 76190 9938
rect 76242 9886 76244 9938
rect 76076 9156 76132 9166
rect 76188 9156 76244 9886
rect 76300 9602 76356 9614
rect 76300 9550 76302 9602
rect 76354 9550 76356 9602
rect 76300 9268 76356 9550
rect 76300 9202 76356 9212
rect 76076 9154 76244 9156
rect 76076 9102 76078 9154
rect 76130 9102 76244 9154
rect 76076 9100 76244 9102
rect 76076 9090 76132 9100
rect 76412 9044 76468 13134
rect 77084 13188 77140 13580
rect 77084 13122 77140 13132
rect 77196 13524 77252 13534
rect 76524 13076 76580 13086
rect 76524 12404 76580 13020
rect 76636 12964 76692 12974
rect 76636 12870 76692 12908
rect 77084 12852 77140 12862
rect 77084 12404 77140 12796
rect 76524 12402 76916 12404
rect 76524 12350 76526 12402
rect 76578 12350 76916 12402
rect 76524 12348 76916 12350
rect 76524 12338 76580 12348
rect 76860 10834 76916 12348
rect 77084 12272 77140 12348
rect 77196 12738 77252 13468
rect 77196 12686 77198 12738
rect 77250 12686 77252 12738
rect 77196 12292 77252 12686
rect 77196 12180 77252 12236
rect 77084 12124 77252 12180
rect 76860 10782 76862 10834
rect 76914 10782 76916 10834
rect 76524 9716 76580 9726
rect 76524 9714 76804 9716
rect 76524 9662 76526 9714
rect 76578 9662 76804 9714
rect 76524 9660 76804 9662
rect 76524 9650 76580 9660
rect 76300 8988 76468 9044
rect 75964 8876 76244 8932
rect 75852 8306 75908 8316
rect 76188 8148 76244 8876
rect 75964 8146 76244 8148
rect 75964 8094 76190 8146
rect 76242 8094 76244 8146
rect 75964 8092 76244 8094
rect 75740 8034 75796 8046
rect 75740 7982 75742 8034
rect 75794 7982 75796 8034
rect 75740 7812 75796 7982
rect 75740 7746 75796 7756
rect 75404 7250 75572 7252
rect 75404 7198 75406 7250
rect 75458 7198 75572 7250
rect 75404 7196 75572 7198
rect 75404 7186 75460 7196
rect 75516 6578 75572 7196
rect 75628 7186 75684 7196
rect 75516 6526 75518 6578
rect 75570 6526 75572 6578
rect 75404 6132 75460 6142
rect 75404 5906 75460 6076
rect 75404 5854 75406 5906
rect 75458 5854 75460 5906
rect 75404 5842 75460 5854
rect 75516 5908 75572 6526
rect 75964 6580 76020 8092
rect 76188 8082 76244 8092
rect 76300 7588 76356 8988
rect 76524 8148 76580 8158
rect 76524 8054 76580 8092
rect 75964 6514 76020 6524
rect 76076 7532 76356 7588
rect 76524 7812 76580 7822
rect 76524 7588 76580 7756
rect 76524 7586 76692 7588
rect 76524 7534 76526 7586
rect 76578 7534 76692 7586
rect 76524 7532 76692 7534
rect 75292 5628 75460 5684
rect 75404 5348 75460 5628
rect 75292 5236 75348 5246
rect 75292 5142 75348 5180
rect 75180 5058 75236 5068
rect 74956 4274 75012 4284
rect 75404 4338 75460 5292
rect 75516 5124 75572 5852
rect 75628 5348 75684 5358
rect 75628 5234 75684 5292
rect 75628 5182 75630 5234
rect 75682 5182 75684 5234
rect 75628 5170 75684 5182
rect 75516 5058 75572 5068
rect 76076 5012 76132 7532
rect 76524 7522 76580 7532
rect 76412 7476 76468 7486
rect 76188 7474 76468 7476
rect 76188 7422 76414 7474
rect 76466 7422 76468 7474
rect 76188 7420 76468 7422
rect 76188 6804 76244 7420
rect 76412 7410 76468 7420
rect 76524 7364 76580 7374
rect 76188 5794 76244 6748
rect 76412 7028 76468 7038
rect 76412 6466 76468 6972
rect 76524 6802 76580 7308
rect 76524 6750 76526 6802
rect 76578 6750 76580 6802
rect 76524 6738 76580 6750
rect 76636 6692 76692 7532
rect 76636 6626 76692 6636
rect 76412 6414 76414 6466
rect 76466 6414 76468 6466
rect 76412 6402 76468 6414
rect 76524 6580 76580 6590
rect 76524 5906 76580 6524
rect 76524 5854 76526 5906
rect 76578 5854 76580 5906
rect 76524 5842 76580 5854
rect 76188 5742 76190 5794
rect 76242 5742 76244 5794
rect 76188 5236 76244 5742
rect 76188 5170 76244 5180
rect 76188 5012 76244 5022
rect 76076 5010 76356 5012
rect 76076 4958 76190 5010
rect 76242 4958 76356 5010
rect 76076 4956 76356 4958
rect 76188 4946 76244 4956
rect 75404 4286 75406 4338
rect 75458 4286 75460 4338
rect 75404 4274 75460 4286
rect 75628 4450 75684 4462
rect 75628 4398 75630 4450
rect 75682 4398 75684 4450
rect 75628 4340 75684 4398
rect 76188 4340 76244 4350
rect 75628 4338 76244 4340
rect 75628 4286 76190 4338
rect 76242 4286 76244 4338
rect 75628 4284 76244 4286
rect 76188 4274 76244 4284
rect 76300 4228 76356 4956
rect 76524 4898 76580 4910
rect 76524 4846 76526 4898
rect 76578 4846 76580 4898
rect 76524 4788 76580 4846
rect 76748 4900 76804 9660
rect 76860 9492 76916 10782
rect 76860 9426 76916 9436
rect 76972 12068 77028 12078
rect 76972 5348 77028 12012
rect 77084 7364 77140 12124
rect 77196 11508 77252 11518
rect 77196 9828 77252 11452
rect 77196 9762 77252 9772
rect 77084 7298 77140 7308
rect 77308 6916 77364 13804
rect 77420 13076 77476 13086
rect 77420 12402 77476 13020
rect 77420 12350 77422 12402
rect 77474 12350 77476 12402
rect 77420 12068 77476 12350
rect 77420 12002 77476 12012
rect 77532 11508 77588 15092
rect 77868 13188 77924 20748
rect 78652 20188 78708 115838
rect 80220 116116 80276 116126
rect 78876 23940 78932 23950
rect 78652 20132 78820 20188
rect 78204 18564 78260 18574
rect 78204 13634 78260 18508
rect 78204 13582 78206 13634
rect 78258 13582 78260 13634
rect 77868 13132 78036 13188
rect 77756 12740 77812 12750
rect 77420 11452 77532 11508
rect 77420 9044 77476 11452
rect 77532 11442 77588 11452
rect 77644 12738 77812 12740
rect 77644 12686 77758 12738
rect 77810 12686 77812 12738
rect 77644 12684 77812 12686
rect 77532 9602 77588 9614
rect 77532 9550 77534 9602
rect 77586 9550 77588 9602
rect 77532 9268 77588 9550
rect 77532 9202 77588 9212
rect 77420 8988 77588 9044
rect 77420 8820 77476 8830
rect 77420 8258 77476 8764
rect 77420 8206 77422 8258
rect 77474 8206 77476 8258
rect 77420 8194 77476 8206
rect 77532 7924 77588 8988
rect 77644 8260 77700 12684
rect 77756 12674 77812 12684
rect 77980 12628 78036 13132
rect 77868 12572 78036 12628
rect 77756 9828 77812 9838
rect 77756 9734 77812 9772
rect 77868 8484 77924 12572
rect 77980 12404 78036 12414
rect 77980 12310 78036 12348
rect 78204 12068 78260 13582
rect 78764 13524 78820 20132
rect 78876 13636 78932 23884
rect 79436 23604 79492 23614
rect 78876 13570 78932 13580
rect 79100 13636 79156 13646
rect 79100 13542 79156 13580
rect 78764 13458 78820 13468
rect 79212 13186 79268 13198
rect 79212 13134 79214 13186
rect 79266 13134 79268 13186
rect 78540 12738 78596 12750
rect 78540 12686 78542 12738
rect 78594 12686 78596 12738
rect 78540 12516 78596 12686
rect 78540 12450 78596 12460
rect 79100 12738 79156 12750
rect 79100 12686 79102 12738
rect 79154 12686 79156 12738
rect 78540 12068 78596 12078
rect 78204 12066 78596 12068
rect 78204 12014 78542 12066
rect 78594 12014 78596 12066
rect 78204 12012 78596 12014
rect 78316 11844 78372 11854
rect 78092 11508 78148 11518
rect 78092 11414 78148 11452
rect 78204 11396 78260 11406
rect 78204 8932 78260 11340
rect 78204 8800 78260 8876
rect 78316 11060 78372 11788
rect 78540 11508 78596 12012
rect 79100 11844 79156 12686
rect 79212 12402 79268 13134
rect 79212 12350 79214 12402
rect 79266 12350 79268 12402
rect 79212 12338 79268 12350
rect 79436 12740 79492 23548
rect 79772 13634 79828 13646
rect 79772 13582 79774 13634
rect 79826 13582 79828 13634
rect 79100 11778 79156 11788
rect 79212 12180 79268 12190
rect 78540 11442 78596 11452
rect 78428 11396 78484 11406
rect 78428 11302 78484 11340
rect 78316 8708 78372 11004
rect 78876 11170 78932 11182
rect 78876 11118 78878 11170
rect 78930 11118 78932 11170
rect 78876 10500 78932 11118
rect 78876 10434 78932 10444
rect 79100 10498 79156 10510
rect 79100 10446 79102 10498
rect 79154 10446 79156 10498
rect 78428 10276 78484 10286
rect 78428 9156 78484 10220
rect 79100 10164 79156 10446
rect 78652 10108 79156 10164
rect 78652 9938 78708 10108
rect 79212 10052 79268 12124
rect 78652 9886 78654 9938
rect 78706 9886 78708 9938
rect 78652 9874 78708 9886
rect 78988 9996 79268 10052
rect 79324 11508 79380 11518
rect 78764 9716 78820 9726
rect 78764 9622 78820 9660
rect 78540 9602 78596 9614
rect 78540 9550 78542 9602
rect 78594 9550 78596 9602
rect 78540 9268 78596 9550
rect 78988 9492 79044 9996
rect 79212 9716 79268 9754
rect 79212 9650 79268 9660
rect 78988 9436 79156 9492
rect 78540 9202 78596 9212
rect 78428 9090 78484 9100
rect 78764 8932 78820 8942
rect 78764 8838 78820 8876
rect 78316 8642 78372 8652
rect 78876 8818 78932 8830
rect 78876 8766 78878 8818
rect 78930 8766 78932 8818
rect 78876 8484 78932 8766
rect 77868 8428 78372 8484
rect 77644 8204 78036 8260
rect 77644 8036 77700 8046
rect 77644 8034 77924 8036
rect 77644 7982 77646 8034
rect 77698 7982 77924 8034
rect 77644 7980 77924 7982
rect 77644 7970 77700 7980
rect 77532 7858 77588 7868
rect 77756 7812 77812 7822
rect 77644 7476 77700 7486
rect 77308 6850 77364 6860
rect 77532 7252 77588 7262
rect 77532 6804 77588 7196
rect 77532 6710 77588 6748
rect 77308 6692 77364 6702
rect 77308 6598 77364 6636
rect 77420 6468 77476 6478
rect 77420 6374 77476 6412
rect 77644 6018 77700 7420
rect 77756 6914 77812 7756
rect 77756 6862 77758 6914
rect 77810 6862 77812 6914
rect 77756 6580 77812 6862
rect 77756 6514 77812 6524
rect 77756 6244 77812 6254
rect 77756 6130 77812 6188
rect 77756 6078 77758 6130
rect 77810 6078 77812 6130
rect 77756 6066 77812 6078
rect 77644 5966 77646 6018
rect 77698 5966 77700 6018
rect 77644 5954 77700 5966
rect 76972 5282 77028 5292
rect 77084 5794 77140 5806
rect 77084 5742 77086 5794
rect 77138 5742 77140 5794
rect 77084 5012 77140 5742
rect 77644 5124 77700 5134
rect 77644 5030 77700 5068
rect 77084 4946 77140 4956
rect 76748 4834 76804 4844
rect 77420 4898 77476 4910
rect 77420 4846 77422 4898
rect 77474 4846 77476 4898
rect 76524 4722 76580 4732
rect 77308 4788 77364 4798
rect 76300 4004 76356 4172
rect 76300 3938 76356 3948
rect 76524 4564 76580 4574
rect 74844 3826 74900 3836
rect 75964 3780 76020 3790
rect 75180 3444 75236 3482
rect 75180 3378 75236 3388
rect 74732 2482 74788 2492
rect 74284 1708 74452 1764
rect 74284 800 74340 1708
rect 75964 800 76020 3724
rect 76524 3666 76580 4508
rect 76860 4226 76916 4238
rect 76860 4174 76862 4226
rect 76914 4174 76916 4226
rect 76860 3780 76916 4174
rect 76860 3714 76916 3724
rect 76972 3892 77028 3902
rect 76972 3778 77028 3836
rect 76972 3726 76974 3778
rect 77026 3726 77028 3778
rect 76972 3714 77028 3726
rect 76524 3614 76526 3666
rect 76578 3614 76580 3666
rect 76524 3602 76580 3614
rect 77084 3668 77140 3678
rect 77084 3574 77140 3612
rect 77308 3554 77364 4732
rect 77420 4676 77476 4846
rect 77420 4610 77476 4620
rect 77532 4898 77588 4910
rect 77532 4846 77534 4898
rect 77586 4846 77588 4898
rect 77532 3668 77588 4846
rect 77532 3602 77588 3612
rect 77308 3502 77310 3554
rect 77362 3502 77364 3554
rect 77308 3490 77364 3502
rect 77868 3554 77924 7980
rect 77980 6356 78036 8204
rect 78204 8146 78260 8158
rect 78204 8094 78206 8146
rect 78258 8094 78260 8146
rect 78204 7252 78260 8094
rect 78316 7252 78372 8428
rect 78764 8428 78932 8484
rect 78540 8372 78596 8382
rect 78540 8278 78596 8316
rect 78428 8146 78484 8158
rect 78428 8094 78430 8146
rect 78482 8094 78484 8146
rect 78428 7812 78484 8094
rect 78428 7746 78484 7756
rect 78540 8148 78596 8158
rect 78540 8036 78596 8092
rect 78764 8036 78820 8428
rect 78988 8260 79044 8270
rect 78988 8166 79044 8204
rect 78540 7980 78820 8036
rect 78540 7474 78596 7980
rect 78540 7422 78542 7474
rect 78594 7422 78596 7474
rect 78540 7410 78596 7422
rect 78876 7924 78932 7934
rect 78316 7196 78596 7252
rect 78204 7186 78260 7196
rect 78092 6916 78148 6926
rect 78092 6580 78148 6860
rect 78428 6580 78484 6590
rect 78092 6524 78260 6580
rect 77980 6132 78036 6300
rect 77980 6076 78148 6132
rect 77980 5908 78036 5918
rect 77980 5814 78036 5852
rect 78092 5906 78148 6076
rect 78092 5854 78094 5906
rect 78146 5854 78148 5906
rect 78092 5842 78148 5854
rect 78204 5234 78260 6524
rect 78428 6486 78484 6524
rect 78204 5182 78206 5234
rect 78258 5182 78260 5234
rect 77980 5012 78036 5022
rect 77980 4918 78036 4956
rect 78092 4900 78148 4910
rect 78092 4806 78148 4844
rect 78204 4452 78260 5182
rect 78204 4386 78260 4396
rect 78428 4900 78484 4910
rect 78428 4450 78484 4844
rect 78540 4562 78596 7196
rect 78764 6580 78820 6590
rect 78876 6580 78932 7868
rect 78988 7588 79044 7598
rect 79100 7588 79156 9436
rect 79324 8146 79380 11452
rect 79436 11506 79492 12684
rect 79436 11454 79438 11506
rect 79490 11454 79492 11506
rect 79436 11442 79492 11454
rect 79548 13186 79604 13198
rect 79548 13134 79550 13186
rect 79602 13134 79604 13186
rect 79324 8094 79326 8146
rect 79378 8094 79380 8146
rect 79212 8034 79268 8046
rect 79212 7982 79214 8034
rect 79266 7982 79268 8034
rect 79212 7924 79268 7982
rect 79212 7858 79268 7868
rect 78988 7586 79156 7588
rect 78988 7534 78990 7586
rect 79042 7534 79156 7586
rect 78988 7532 79156 7534
rect 78988 7522 79044 7532
rect 78764 6578 78932 6580
rect 78764 6526 78766 6578
rect 78818 6526 78932 6578
rect 78764 6524 78932 6526
rect 78764 6514 78820 6524
rect 78876 6244 78932 6254
rect 78876 5906 78932 6188
rect 79100 6020 79156 6030
rect 79100 6018 79268 6020
rect 79100 5966 79102 6018
rect 79154 5966 79268 6018
rect 79100 5964 79268 5966
rect 79100 5954 79156 5964
rect 78876 5854 78878 5906
rect 78930 5854 78932 5906
rect 78876 5842 78932 5854
rect 78988 5908 79044 5918
rect 78652 5236 78708 5246
rect 78652 5142 78708 5180
rect 78540 4510 78542 4562
rect 78594 4510 78596 4562
rect 78540 4498 78596 4510
rect 78652 5012 78708 5022
rect 78988 5012 79044 5852
rect 79100 5012 79156 5022
rect 78988 5010 79156 5012
rect 78988 4958 79102 5010
rect 79154 4958 79156 5010
rect 78988 4956 79156 4958
rect 78652 4788 78708 4956
rect 79100 4946 79156 4956
rect 78652 4562 78708 4732
rect 78652 4510 78654 4562
rect 78706 4510 78708 4562
rect 78652 4498 78708 4510
rect 78428 4398 78430 4450
rect 78482 4398 78484 4450
rect 78428 4386 78484 4398
rect 79212 4340 79268 5964
rect 79324 4900 79380 8094
rect 79436 6916 79492 6926
rect 79436 5010 79492 6860
rect 79548 6692 79604 13134
rect 79772 13186 79828 13582
rect 80220 13524 80276 116060
rect 80780 23044 80836 23054
rect 80220 13458 80276 13468
rect 80556 16884 80612 16894
rect 80556 13636 80612 16828
rect 80668 13636 80724 13646
rect 80556 13634 80724 13636
rect 80556 13582 80670 13634
rect 80722 13582 80724 13634
rect 80556 13580 80724 13582
rect 79772 13134 79774 13186
rect 79826 13134 79828 13186
rect 79772 13122 79828 13134
rect 79660 12852 79716 12862
rect 79660 12758 79716 12796
rect 79884 12852 79940 12862
rect 79660 12066 79716 12078
rect 79660 12014 79662 12066
rect 79714 12014 79716 12066
rect 79660 11844 79716 12014
rect 79660 11778 79716 11788
rect 79772 10610 79828 10622
rect 79772 10558 79774 10610
rect 79826 10558 79828 10610
rect 79772 10500 79828 10558
rect 79772 10434 79828 10444
rect 79660 9602 79716 9614
rect 79660 9550 79662 9602
rect 79714 9550 79716 9602
rect 79660 9492 79716 9550
rect 79660 9426 79716 9436
rect 79660 9268 79716 9278
rect 79660 9174 79716 9212
rect 79884 8372 79940 12796
rect 79996 12740 80052 12750
rect 80556 12740 80612 13580
rect 80668 13570 80724 13580
rect 79996 12738 80612 12740
rect 79996 12686 79998 12738
rect 80050 12686 80612 12738
rect 79996 12684 80612 12686
rect 79996 12674 80052 12684
rect 79772 8316 79940 8372
rect 79996 12516 80052 12526
rect 79772 7700 79828 8316
rect 79772 6916 79828 7644
rect 79884 8148 79940 8158
rect 79884 7588 79940 8092
rect 79884 7522 79940 7532
rect 79772 6850 79828 6860
rect 79660 6692 79716 6702
rect 79548 6690 79716 6692
rect 79548 6638 79662 6690
rect 79714 6638 79716 6690
rect 79548 6636 79716 6638
rect 79996 6692 80052 12460
rect 80108 12068 80164 12078
rect 80108 11974 80164 12012
rect 80108 9604 80164 9614
rect 80108 9510 80164 9548
rect 80108 8932 80164 8942
rect 80108 8838 80164 8876
rect 80108 8596 80164 8606
rect 80108 7698 80164 8540
rect 80108 7646 80110 7698
rect 80162 7646 80164 7698
rect 80108 7634 80164 7646
rect 80220 8034 80276 8046
rect 80220 7982 80222 8034
rect 80274 7982 80276 8034
rect 79996 6636 80164 6692
rect 79660 5796 79716 6636
rect 79772 6580 79828 6590
rect 79772 6486 79828 6524
rect 79996 6466 80052 6478
rect 79996 6414 79998 6466
rect 80050 6414 80052 6466
rect 79884 6356 79940 6366
rect 79884 6130 79940 6300
rect 79884 6078 79886 6130
rect 79938 6078 79940 6130
rect 79884 6066 79940 6078
rect 79996 6020 80052 6414
rect 80108 6132 80164 6636
rect 80108 6066 80164 6076
rect 79996 5954 80052 5964
rect 79660 5740 80052 5796
rect 79996 5348 80052 5740
rect 80220 5684 80276 7982
rect 80332 5908 80388 12684
rect 80556 12516 80612 12526
rect 80556 12402 80612 12460
rect 80556 12350 80558 12402
rect 80610 12350 80612 12402
rect 80556 12338 80612 12350
rect 80444 10500 80500 10510
rect 80444 10498 80612 10500
rect 80444 10446 80446 10498
rect 80498 10446 80612 10498
rect 80444 10444 80612 10446
rect 80444 10434 80500 10444
rect 80444 9268 80500 9278
rect 80444 8484 80500 9212
rect 80444 8418 80500 8428
rect 80556 9266 80612 10444
rect 80556 9214 80558 9266
rect 80610 9214 80612 9266
rect 80556 8820 80612 9214
rect 80556 8148 80612 8764
rect 80668 9602 80724 9614
rect 80668 9550 80670 9602
rect 80722 9550 80724 9602
rect 80668 8596 80724 9550
rect 80780 9268 80836 22988
rect 81116 23044 81172 116396
rect 81228 116386 81284 116396
rect 81900 116386 81956 116396
rect 81276 116060 81540 116070
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81276 115994 81540 116004
rect 82908 115892 82964 119200
rect 84476 117908 84532 119200
rect 84476 117852 84980 117908
rect 84924 116562 84980 117852
rect 84924 116510 84926 116562
rect 84978 116510 84980 116562
rect 84924 116498 84980 116510
rect 85932 116450 85988 116462
rect 85932 116398 85934 116450
rect 85986 116398 85988 116450
rect 85932 116116 85988 116398
rect 85932 116050 85988 116060
rect 86380 116226 86436 116238
rect 86380 116174 86382 116226
rect 86434 116174 86436 116226
rect 86380 116116 86436 116174
rect 86380 116050 86436 116060
rect 82908 115826 82964 115836
rect 83804 115892 83860 115902
rect 82572 115778 82628 115790
rect 82572 115726 82574 115778
rect 82626 115726 82628 115778
rect 82236 115666 82292 115678
rect 82236 115614 82238 115666
rect 82290 115614 82292 115666
rect 81676 115556 81732 115566
rect 81676 115462 81732 115500
rect 82236 115556 82292 115614
rect 82572 115668 82628 115726
rect 83132 115668 83188 115678
rect 82572 115666 83188 115668
rect 82572 115614 83134 115666
rect 83186 115614 83188 115666
rect 82572 115612 83188 115614
rect 83132 115602 83188 115612
rect 82236 114884 82292 115500
rect 83804 115554 83860 115836
rect 83804 115502 83806 115554
rect 83858 115502 83860 115554
rect 83804 115490 83860 115502
rect 87276 115666 87332 115678
rect 87276 115614 87278 115666
rect 87330 115614 87332 115666
rect 82236 114818 82292 114828
rect 86716 114884 86772 114894
rect 86716 114790 86772 114828
rect 87276 114770 87332 115614
rect 87612 115556 87668 119200
rect 89180 117908 89236 119200
rect 89180 117852 89684 117908
rect 89628 116562 89684 117852
rect 92316 116676 92372 119200
rect 92316 116610 92372 116620
rect 93212 116676 93268 116686
rect 89628 116510 89630 116562
rect 89682 116510 89684 116562
rect 89628 116498 89684 116510
rect 93212 116562 93268 116620
rect 93212 116510 93214 116562
rect 93266 116510 93268 116562
rect 93212 116498 93268 116510
rect 90636 116450 90692 116462
rect 92540 116452 92596 116462
rect 90636 116398 90638 116450
rect 90690 116398 90692 116450
rect 90636 116228 90692 116398
rect 92316 116450 92596 116452
rect 92316 116398 92542 116450
rect 92594 116398 92596 116450
rect 92316 116396 92596 116398
rect 90636 116162 90692 116172
rect 91084 116228 91140 116238
rect 91084 116134 91140 116172
rect 90860 116116 90916 116126
rect 87948 115556 88004 115566
rect 87612 115554 88004 115556
rect 87612 115502 87950 115554
rect 88002 115502 88004 115554
rect 87612 115500 88004 115502
rect 87948 115490 88004 115500
rect 87612 114884 87668 114894
rect 87612 114790 87668 114828
rect 87276 114718 87278 114770
rect 87330 114718 87332 114770
rect 87276 114706 87332 114718
rect 81276 114492 81540 114502
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81276 114426 81540 114436
rect 81276 112924 81540 112934
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81276 112858 81540 112868
rect 81276 111356 81540 111366
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81276 111290 81540 111300
rect 81276 109788 81540 109798
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81276 109722 81540 109732
rect 81276 108220 81540 108230
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81276 108154 81540 108164
rect 81276 106652 81540 106662
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81276 106586 81540 106596
rect 81276 105084 81540 105094
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81276 105018 81540 105028
rect 81276 103516 81540 103526
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81276 103450 81540 103460
rect 81276 101948 81540 101958
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81276 101882 81540 101892
rect 81276 100380 81540 100390
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81276 100314 81540 100324
rect 81276 98812 81540 98822
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81276 98746 81540 98756
rect 81276 97244 81540 97254
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81276 97178 81540 97188
rect 81276 95676 81540 95686
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81276 95610 81540 95620
rect 81276 94108 81540 94118
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81276 94042 81540 94052
rect 81276 92540 81540 92550
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81276 92474 81540 92484
rect 81276 90972 81540 90982
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81276 90906 81540 90916
rect 81276 89404 81540 89414
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81276 89338 81540 89348
rect 81276 87836 81540 87846
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81276 87770 81540 87780
rect 81276 86268 81540 86278
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81276 86202 81540 86212
rect 81276 84700 81540 84710
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81276 84634 81540 84644
rect 81276 83132 81540 83142
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81276 83066 81540 83076
rect 81276 81564 81540 81574
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81276 81498 81540 81508
rect 81276 79996 81540 80006
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81276 79930 81540 79940
rect 81276 78428 81540 78438
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81276 78362 81540 78372
rect 81276 76860 81540 76870
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81276 76794 81540 76804
rect 81276 75292 81540 75302
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81276 75226 81540 75236
rect 81276 73724 81540 73734
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81276 73658 81540 73668
rect 81276 72156 81540 72166
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81276 72090 81540 72100
rect 81276 70588 81540 70598
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81276 70522 81540 70532
rect 81276 69020 81540 69030
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81276 68954 81540 68964
rect 81276 67452 81540 67462
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81276 67386 81540 67396
rect 81276 65884 81540 65894
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81276 65818 81540 65828
rect 81276 64316 81540 64326
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81276 64250 81540 64260
rect 81276 62748 81540 62758
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81276 62682 81540 62692
rect 81276 61180 81540 61190
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81276 61114 81540 61124
rect 81276 59612 81540 59622
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81276 59546 81540 59556
rect 81276 58044 81540 58054
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81276 57978 81540 57988
rect 81276 56476 81540 56486
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81276 56410 81540 56420
rect 81276 54908 81540 54918
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81276 54842 81540 54852
rect 81276 53340 81540 53350
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81276 53274 81540 53284
rect 81276 51772 81540 51782
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81276 51706 81540 51716
rect 81276 50204 81540 50214
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81276 50138 81540 50148
rect 81276 48636 81540 48646
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81276 48570 81540 48580
rect 81276 47068 81540 47078
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81276 47002 81540 47012
rect 81276 45500 81540 45510
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81276 45434 81540 45444
rect 81276 43932 81540 43942
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81276 43866 81540 43876
rect 81276 42364 81540 42374
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81276 42298 81540 42308
rect 81276 40796 81540 40806
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81276 40730 81540 40740
rect 81276 39228 81540 39238
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81276 39162 81540 39172
rect 81276 37660 81540 37670
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81276 37594 81540 37604
rect 81276 36092 81540 36102
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81276 36026 81540 36036
rect 81276 34524 81540 34534
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81276 34458 81540 34468
rect 81276 32956 81540 32966
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81276 32890 81540 32900
rect 81276 31388 81540 31398
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81276 31322 81540 31332
rect 81276 29820 81540 29830
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81276 29754 81540 29764
rect 81276 28252 81540 28262
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81276 28186 81540 28196
rect 81276 26684 81540 26694
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81276 26618 81540 26628
rect 90860 25620 90916 116060
rect 92316 115890 92372 116396
rect 92540 116386 92596 116396
rect 92316 115838 92318 115890
rect 92370 115838 92372 115890
rect 92316 115826 92372 115838
rect 93884 115780 93940 119200
rect 96636 116844 96900 116854
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96636 116778 96900 116788
rect 97020 116564 97076 119200
rect 97020 116498 97076 116508
rect 97916 116564 97972 116574
rect 97916 116470 97972 116508
rect 98588 116564 98644 119200
rect 101724 116676 101780 119200
rect 101724 116610 101780 116620
rect 102508 116676 102564 116686
rect 98588 116498 98644 116508
rect 100044 116564 100100 116574
rect 100044 116470 100100 116508
rect 102508 116562 102564 116620
rect 102508 116510 102510 116562
rect 102562 116510 102564 116562
rect 102508 116498 102564 116510
rect 103292 116564 103348 119200
rect 103292 116498 103348 116508
rect 104188 116564 104244 116574
rect 104188 116470 104244 116508
rect 106428 116564 106484 119200
rect 106428 116498 106484 116508
rect 97244 116450 97300 116462
rect 97244 116398 97246 116450
rect 97298 116398 97300 116450
rect 97244 115890 97300 116398
rect 97244 115838 97246 115890
rect 97298 115838 97300 115890
rect 97244 115826 97300 115838
rect 101052 116450 101108 116462
rect 101052 116398 101054 116450
rect 101106 116398 101108 116450
rect 93884 115714 93940 115724
rect 94444 115780 94500 115790
rect 94444 115686 94500 115724
rect 91420 115668 91476 115678
rect 91420 115554 91476 115612
rect 91980 115668 92036 115678
rect 91980 115574 92036 115612
rect 95340 115666 95396 115678
rect 95340 115614 95342 115666
rect 95394 115614 95396 115666
rect 91420 115502 91422 115554
rect 91474 115502 91476 115554
rect 91420 114884 91476 115502
rect 95340 115556 95396 115614
rect 96460 115668 96516 115678
rect 96460 115574 96516 115612
rect 97580 115668 97636 115678
rect 97580 115574 97636 115612
rect 100828 115668 100884 115678
rect 100828 115574 100884 115612
rect 95340 115490 95396 115500
rect 95900 115556 95956 115566
rect 95900 115462 95956 115500
rect 97468 115556 97524 115566
rect 96636 115276 96900 115286
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96636 115210 96900 115220
rect 91420 114818 91476 114828
rect 96636 113708 96900 113718
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96636 113642 96900 113652
rect 96636 112140 96900 112150
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96636 112074 96900 112084
rect 96636 110572 96900 110582
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96636 110506 96900 110516
rect 96636 109004 96900 109014
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96636 108938 96900 108948
rect 96636 107436 96900 107446
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96636 107370 96900 107380
rect 96636 105868 96900 105878
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96636 105802 96900 105812
rect 96636 104300 96900 104310
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96636 104234 96900 104244
rect 96636 102732 96900 102742
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96636 102666 96900 102676
rect 96636 101164 96900 101174
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96636 101098 96900 101108
rect 96636 99596 96900 99606
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96636 99530 96900 99540
rect 96636 98028 96900 98038
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96636 97962 96900 97972
rect 96636 96460 96900 96470
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96636 96394 96900 96404
rect 96636 94892 96900 94902
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96636 94826 96900 94836
rect 96636 93324 96900 93334
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96636 93258 96900 93268
rect 96636 91756 96900 91766
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96636 91690 96900 91700
rect 96636 90188 96900 90198
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96636 90122 96900 90132
rect 96636 88620 96900 88630
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96636 88554 96900 88564
rect 96636 87052 96900 87062
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96636 86986 96900 86996
rect 96636 85484 96900 85494
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96636 85418 96900 85428
rect 96636 83916 96900 83926
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96636 83850 96900 83860
rect 96636 82348 96900 82358
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96636 82282 96900 82292
rect 96636 80780 96900 80790
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96636 80714 96900 80724
rect 96636 79212 96900 79222
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96636 79146 96900 79156
rect 96636 77644 96900 77654
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96636 77578 96900 77588
rect 96636 76076 96900 76086
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96636 76010 96900 76020
rect 96636 74508 96900 74518
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96636 74442 96900 74452
rect 96636 72940 96900 72950
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96636 72874 96900 72884
rect 96636 71372 96900 71382
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96636 71306 96900 71316
rect 96636 69804 96900 69814
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96636 69738 96900 69748
rect 96636 68236 96900 68246
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96636 68170 96900 68180
rect 96636 66668 96900 66678
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96636 66602 96900 66612
rect 96636 65100 96900 65110
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96636 65034 96900 65044
rect 96636 63532 96900 63542
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96636 63466 96900 63476
rect 96636 61964 96900 61974
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96636 61898 96900 61908
rect 96636 60396 96900 60406
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96636 60330 96900 60340
rect 96636 58828 96900 58838
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96636 58762 96900 58772
rect 96636 57260 96900 57270
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96636 57194 96900 57204
rect 96636 55692 96900 55702
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96636 55626 96900 55636
rect 96636 54124 96900 54134
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96636 54058 96900 54068
rect 96636 52556 96900 52566
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96636 52490 96900 52500
rect 96636 50988 96900 50998
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96636 50922 96900 50932
rect 96636 49420 96900 49430
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96636 49354 96900 49364
rect 96636 47852 96900 47862
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96636 47786 96900 47796
rect 96636 46284 96900 46294
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96636 46218 96900 46228
rect 96636 44716 96900 44726
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96636 44650 96900 44660
rect 96636 43148 96900 43158
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96636 43082 96900 43092
rect 96636 41580 96900 41590
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96636 41514 96900 41524
rect 96636 40012 96900 40022
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96636 39946 96900 39956
rect 96636 38444 96900 38454
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96636 38378 96900 38388
rect 96636 36876 96900 36886
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96636 36810 96900 36820
rect 96636 35308 96900 35318
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96636 35242 96900 35252
rect 96636 33740 96900 33750
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96636 33674 96900 33684
rect 96636 32172 96900 32182
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96636 32106 96900 32116
rect 96636 30604 96900 30614
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96636 30538 96900 30548
rect 96636 29036 96900 29046
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96636 28970 96900 28980
rect 96636 27468 96900 27478
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96636 27402 96900 27412
rect 97468 27300 97524 115500
rect 101052 115444 101108 116398
rect 101724 116450 101780 116462
rect 101724 116398 101726 116450
rect 101778 116398 101780 116450
rect 101724 115890 101780 116398
rect 104972 116450 105028 116462
rect 104972 116398 104974 116450
rect 105026 116398 105028 116450
rect 104972 116228 105028 116398
rect 106316 116452 106372 116462
rect 104972 116162 105028 116172
rect 105420 116228 105476 116238
rect 105420 116134 105476 116172
rect 106092 116228 106148 116238
rect 101724 115838 101726 115890
rect 101778 115838 101780 115890
rect 101724 115826 101780 115838
rect 101388 115668 101444 115678
rect 101388 115574 101444 115612
rect 105420 115668 105476 115678
rect 105420 115574 105476 115612
rect 105980 115668 106036 115678
rect 105980 115574 106036 115612
rect 102172 115554 102228 115566
rect 102172 115502 102174 115554
rect 102226 115502 102228 115554
rect 102172 115444 102228 115502
rect 101052 115388 102228 115444
rect 97468 27234 97524 27244
rect 98364 27300 98420 27310
rect 96636 25900 96900 25910
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96636 25834 96900 25844
rect 90860 25554 90916 25564
rect 91532 25620 91588 25630
rect 81276 25116 81540 25126
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81276 25050 81540 25060
rect 81276 23548 81540 23558
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81276 23482 81540 23492
rect 81116 22978 81172 22988
rect 82012 22260 82068 22270
rect 81276 21980 81540 21990
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81276 21914 81540 21924
rect 81276 20412 81540 20422
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81276 20346 81540 20356
rect 81004 19460 81060 19470
rect 80892 12738 80948 12750
rect 80892 12686 80894 12738
rect 80946 12686 80948 12738
rect 80892 11844 80948 12686
rect 80892 11778 80948 11788
rect 81004 10052 81060 19404
rect 81276 18844 81540 18854
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81276 18778 81540 18788
rect 81276 17276 81540 17286
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81276 17210 81540 17220
rect 81276 15708 81540 15718
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81276 15642 81540 15652
rect 81276 14140 81540 14150
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81276 14074 81540 14084
rect 82012 12852 82068 22204
rect 84812 20692 84868 20702
rect 82348 18676 82404 18686
rect 80780 9202 80836 9212
rect 80892 9996 81060 10052
rect 81116 12740 81172 12750
rect 80668 8530 80724 8540
rect 80780 8932 80836 8942
rect 80556 8082 80612 8092
rect 80668 8372 80724 8382
rect 80668 8258 80724 8316
rect 80668 8206 80670 8258
rect 80722 8206 80724 8258
rect 80668 6802 80724 8206
rect 80780 7700 80836 8876
rect 80892 8484 80948 9996
rect 81004 9828 81060 9838
rect 81004 9734 81060 9772
rect 81004 9492 81060 9502
rect 81004 9156 81060 9436
rect 81116 9268 81172 12684
rect 81452 12740 81508 12778
rect 81452 12674 81508 12684
rect 81276 12572 81540 12582
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81276 12506 81540 12516
rect 81676 12404 81732 12414
rect 81676 12310 81732 12348
rect 82012 12404 82068 12796
rect 82012 12338 82068 12348
rect 82124 12964 82180 12974
rect 81340 12066 81396 12078
rect 81340 12014 81342 12066
rect 81394 12014 81396 12066
rect 81340 11844 81396 12014
rect 81340 11778 81396 11788
rect 82124 11732 82180 12908
rect 82236 12068 82292 12078
rect 82348 12068 82404 18620
rect 83020 13524 83076 13534
rect 83020 13076 83076 13468
rect 83020 12944 83076 13020
rect 82684 12738 82740 12750
rect 82684 12686 82686 12738
rect 82738 12686 82740 12738
rect 82572 12404 82628 12414
rect 82572 12310 82628 12348
rect 82292 12012 82404 12068
rect 82236 11974 82292 12012
rect 82012 11676 82180 11732
rect 82348 11844 82404 11854
rect 81564 11284 81620 11294
rect 81564 11282 81732 11284
rect 81564 11230 81566 11282
rect 81618 11230 81732 11282
rect 81564 11228 81732 11230
rect 81564 11218 81620 11228
rect 81276 11004 81540 11014
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81276 10938 81540 10948
rect 81228 10500 81284 10510
rect 81228 10406 81284 10444
rect 81676 10052 81732 11228
rect 81676 9986 81732 9996
rect 81788 10610 81844 10622
rect 81788 10558 81790 10610
rect 81842 10558 81844 10610
rect 81452 9828 81508 9838
rect 81452 9734 81508 9772
rect 81788 9828 81844 10558
rect 81788 9762 81844 9772
rect 81276 9436 81540 9446
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81276 9370 81540 9380
rect 81564 9268 81620 9278
rect 81116 9212 81564 9268
rect 82012 9268 82068 11676
rect 82124 11508 82180 11518
rect 82124 10834 82180 11452
rect 82124 10782 82126 10834
rect 82178 10782 82180 10834
rect 82124 10770 82180 10782
rect 82236 11394 82292 11406
rect 82236 11342 82238 11394
rect 82290 11342 82292 11394
rect 82236 10500 82292 11342
rect 82236 10434 82292 10444
rect 82236 9828 82292 9838
rect 82236 9734 82292 9772
rect 82348 9604 82404 11788
rect 82684 10948 82740 12686
rect 83244 12066 83300 12078
rect 83692 12068 83748 12078
rect 84140 12068 84196 12078
rect 83244 12014 83246 12066
rect 83298 12014 83300 12066
rect 83244 11844 83300 12014
rect 83244 11778 83300 11788
rect 83356 12066 83748 12068
rect 83356 12014 83694 12066
rect 83746 12014 83748 12066
rect 83356 12012 83748 12014
rect 82796 11508 82852 11518
rect 82796 11414 82852 11452
rect 82684 10892 82852 10948
rect 82684 10724 82740 10734
rect 82684 10610 82740 10668
rect 82684 10558 82686 10610
rect 82738 10558 82740 10610
rect 82684 10500 82740 10558
rect 82684 10434 82740 10444
rect 82348 9538 82404 9548
rect 82572 9602 82628 9614
rect 82572 9550 82574 9602
rect 82626 9550 82628 9602
rect 82572 9492 82628 9550
rect 82572 9426 82628 9436
rect 82572 9268 82628 9278
rect 82012 9212 82292 9268
rect 81004 9100 81172 9156
rect 81564 9136 81620 9212
rect 80892 8428 81060 8484
rect 80892 8260 80948 8270
rect 80892 8166 80948 8204
rect 80780 7634 80836 7644
rect 81004 7476 81060 8428
rect 81004 7410 81060 7420
rect 81116 8258 81172 9100
rect 82124 9044 82180 9054
rect 82012 9042 82180 9044
rect 82012 8990 82126 9042
rect 82178 8990 82180 9042
rect 82012 8988 82180 8990
rect 81900 8708 81956 8718
rect 81788 8484 81844 8494
rect 81116 8206 81118 8258
rect 81170 8206 81172 8258
rect 81116 7252 81172 8206
rect 81676 8372 81732 8382
rect 81340 8148 81396 8158
rect 81340 8054 81396 8092
rect 81276 7868 81540 7878
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81276 7802 81540 7812
rect 81564 7700 81620 7710
rect 81564 7586 81620 7644
rect 81564 7534 81566 7586
rect 81618 7534 81620 7586
rect 81564 7522 81620 7534
rect 81676 7698 81732 8316
rect 81676 7646 81678 7698
rect 81730 7646 81732 7698
rect 81676 7588 81732 7646
rect 81676 7522 81732 7532
rect 80668 6750 80670 6802
rect 80722 6750 80724 6802
rect 80668 6738 80724 6750
rect 80780 7196 81172 7252
rect 81228 7476 81284 7486
rect 80780 6690 80836 7196
rect 80780 6638 80782 6690
rect 80834 6638 80836 6690
rect 80332 5814 80388 5852
rect 80444 6580 80500 6590
rect 80444 6018 80500 6524
rect 80780 6244 80836 6638
rect 81228 6804 81284 7420
rect 81676 7252 81732 7262
rect 81676 7158 81732 7196
rect 81228 6468 81284 6748
rect 81452 6580 81508 6590
rect 81452 6486 81508 6524
rect 80780 6178 80836 6188
rect 81004 6412 81284 6468
rect 80444 5966 80446 6018
rect 80498 5966 80500 6018
rect 80220 5628 80388 5684
rect 79436 4958 79438 5010
rect 79490 4958 79492 5010
rect 79436 4946 79492 4958
rect 79884 5346 80052 5348
rect 79884 5294 79998 5346
rect 80050 5294 80052 5346
rect 79884 5292 80052 5294
rect 79324 4834 79380 4844
rect 79324 4340 79380 4350
rect 79212 4338 79380 4340
rect 79212 4286 79326 4338
rect 79378 4286 79380 4338
rect 79212 4284 79380 4286
rect 79324 4274 79380 4284
rect 77980 4228 78036 4238
rect 77980 4134 78036 4172
rect 77868 3502 77870 3554
rect 77922 3502 77924 3554
rect 77868 3490 77924 3502
rect 79324 3780 79380 3790
rect 77644 3444 77700 3454
rect 77644 800 77700 3388
rect 78764 3444 78820 3482
rect 78764 3378 78820 3388
rect 79324 800 79380 3724
rect 79884 1652 79940 5292
rect 79996 5282 80052 5292
rect 80220 5012 80276 5022
rect 80220 4918 80276 4956
rect 80108 4900 80164 4910
rect 80108 4806 80164 4844
rect 79996 4226 80052 4238
rect 79996 4174 79998 4226
rect 80050 4174 80052 4226
rect 79996 3780 80052 4174
rect 79996 3714 80052 3724
rect 80332 3554 80388 5628
rect 80444 4004 80500 5966
rect 80668 5908 80724 5918
rect 80668 5814 80724 5852
rect 80892 5796 80948 5806
rect 80892 5346 80948 5740
rect 80892 5294 80894 5346
rect 80946 5294 80948 5346
rect 80892 5282 80948 5294
rect 81004 4564 81060 6412
rect 81276 6300 81540 6310
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81276 6234 81540 6244
rect 81452 6132 81508 6142
rect 81452 6038 81508 6076
rect 81676 6132 81732 6142
rect 81788 6132 81844 8428
rect 81676 6130 81844 6132
rect 81676 6078 81678 6130
rect 81730 6078 81844 6130
rect 81676 6076 81844 6078
rect 81676 6066 81732 6076
rect 81340 6020 81396 6030
rect 81340 5926 81396 5964
rect 81228 5236 81284 5246
rect 81228 5142 81284 5180
rect 81900 5122 81956 8652
rect 82012 8260 82068 8988
rect 82124 8978 82180 8988
rect 82124 8820 82180 8830
rect 82124 8726 82180 8764
rect 82012 8194 82068 8204
rect 82124 8372 82180 8382
rect 82124 7700 82180 8316
rect 81900 5070 81902 5122
rect 81954 5070 81956 5122
rect 81900 5058 81956 5070
rect 82012 7644 82180 7700
rect 81116 5012 81172 5022
rect 81116 4918 81172 4956
rect 81276 4732 81540 4742
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81276 4666 81540 4676
rect 81564 4564 81620 4574
rect 81004 4562 81620 4564
rect 81004 4510 81566 4562
rect 81618 4510 81620 4562
rect 81004 4508 81620 4510
rect 81564 4498 81620 4508
rect 80444 3938 80500 3948
rect 82012 4450 82068 7644
rect 82236 7588 82292 9212
rect 82124 7532 82292 7588
rect 82460 8818 82516 8830
rect 82460 8766 82462 8818
rect 82514 8766 82516 8818
rect 82460 8370 82516 8766
rect 82460 8318 82462 8370
rect 82514 8318 82516 8370
rect 82124 7140 82180 7532
rect 82348 7476 82404 7486
rect 82348 7382 82404 7420
rect 82460 7252 82516 8318
rect 82572 8708 82628 9212
rect 82572 8258 82628 8652
rect 82572 8206 82574 8258
rect 82626 8206 82628 8258
rect 82572 8194 82628 8206
rect 82124 7074 82180 7084
rect 82348 7196 82516 7252
rect 82236 6916 82292 6926
rect 82124 6690 82180 6702
rect 82124 6638 82126 6690
rect 82178 6638 82180 6690
rect 82124 5908 82180 6638
rect 82236 6578 82292 6860
rect 82236 6526 82238 6578
rect 82290 6526 82292 6578
rect 82236 6514 82292 6526
rect 82348 6468 82404 7196
rect 82348 6402 82404 6412
rect 82460 6466 82516 6478
rect 82460 6414 82462 6466
rect 82514 6414 82516 6466
rect 82124 5814 82180 5852
rect 82236 6356 82292 6366
rect 82012 4398 82014 4450
rect 82066 4398 82068 4450
rect 80332 3502 80334 3554
rect 80386 3502 80388 3554
rect 80332 3490 80388 3502
rect 81004 3666 81060 3678
rect 81004 3614 81006 3666
rect 81058 3614 81060 3666
rect 79884 1586 79940 1596
rect 81004 800 81060 3614
rect 81276 3164 81540 3174
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81276 3098 81540 3108
rect 82012 1316 82068 4398
rect 82124 4898 82180 4910
rect 82124 4846 82126 4898
rect 82178 4846 82180 4898
rect 82124 3554 82180 4846
rect 82236 4564 82292 6300
rect 82460 6244 82516 6414
rect 82460 6178 82516 6188
rect 82684 6356 82740 6366
rect 82348 6132 82404 6142
rect 82348 6038 82404 6076
rect 82572 6132 82628 6142
rect 82572 6038 82628 6076
rect 82684 6020 82740 6300
rect 82796 6132 82852 10892
rect 82908 9604 82964 9614
rect 82908 6690 82964 9548
rect 83132 9604 83188 9614
rect 83132 9510 83188 9548
rect 83020 9044 83076 9054
rect 83020 8950 83076 8988
rect 83356 8372 83412 12012
rect 83692 12002 83748 12012
rect 84028 12066 84196 12068
rect 84028 12014 84142 12066
rect 84194 12014 84196 12066
rect 84028 12012 84196 12014
rect 83468 11508 83524 11518
rect 83468 11282 83524 11452
rect 83468 11230 83470 11282
rect 83522 11230 83524 11282
rect 83468 11218 83524 11230
rect 83692 11282 83748 11294
rect 83692 11230 83694 11282
rect 83746 11230 83748 11282
rect 83580 11170 83636 11182
rect 83580 11118 83582 11170
rect 83634 11118 83636 11170
rect 83468 10724 83524 10734
rect 83580 10724 83636 11118
rect 83468 10722 83636 10724
rect 83468 10670 83470 10722
rect 83522 10670 83636 10722
rect 83468 10668 83636 10670
rect 83468 10658 83524 10668
rect 83580 10052 83636 10062
rect 83580 9958 83636 9996
rect 83692 9828 83748 11230
rect 82908 6638 82910 6690
rect 82962 6638 82964 6690
rect 82908 6356 82964 6638
rect 82908 6290 82964 6300
rect 83020 8316 83412 8372
rect 83468 9772 83748 9828
rect 83020 7028 83076 8316
rect 83244 8146 83300 8158
rect 83244 8094 83246 8146
rect 83298 8094 83300 8146
rect 82796 6076 82964 6132
rect 82684 5906 82740 5964
rect 82684 5854 82686 5906
rect 82738 5854 82740 5906
rect 82684 5842 82740 5854
rect 82236 4498 82292 4508
rect 82460 5794 82516 5806
rect 82460 5742 82462 5794
rect 82514 5742 82516 5794
rect 82348 4452 82404 4462
rect 82460 4452 82516 5742
rect 82684 5348 82740 5358
rect 82684 4898 82740 5292
rect 82684 4846 82686 4898
rect 82738 4846 82740 4898
rect 82684 4834 82740 4846
rect 82460 4396 82852 4452
rect 82348 4358 82404 4396
rect 82796 4338 82852 4396
rect 82796 4286 82798 4338
rect 82850 4286 82852 4338
rect 82796 4274 82852 4286
rect 82908 4340 82964 6076
rect 83020 5796 83076 6972
rect 83132 7362 83188 7374
rect 83132 7310 83134 7362
rect 83186 7310 83188 7362
rect 83132 6914 83188 7310
rect 83132 6862 83134 6914
rect 83186 6862 83188 6914
rect 83132 6132 83188 6862
rect 83132 6066 83188 6076
rect 83244 5908 83300 8094
rect 83468 7700 83524 9772
rect 83916 9716 83972 9726
rect 83804 9714 83972 9716
rect 83804 9662 83918 9714
rect 83970 9662 83972 9714
rect 83804 9660 83972 9662
rect 83692 9602 83748 9614
rect 83692 9550 83694 9602
rect 83746 9550 83748 9602
rect 83692 9492 83748 9550
rect 83692 9426 83748 9436
rect 83580 8932 83636 8942
rect 83580 8838 83636 8876
rect 83692 8372 83748 8382
rect 83692 8278 83748 8316
rect 83468 7644 83748 7700
rect 83468 7476 83524 7486
rect 83468 6914 83524 7420
rect 83468 6862 83470 6914
rect 83522 6862 83524 6914
rect 83468 6356 83524 6862
rect 83244 5842 83300 5852
rect 83356 6300 83468 6356
rect 83020 5348 83076 5740
rect 83356 5684 83412 6300
rect 83468 6290 83524 6300
rect 83468 6132 83524 6142
rect 83468 5906 83524 6076
rect 83468 5854 83470 5906
rect 83522 5854 83524 5906
rect 83468 5842 83524 5854
rect 83020 5282 83076 5292
rect 83244 5628 83412 5684
rect 82908 4274 82964 4284
rect 83244 4338 83300 5628
rect 83580 5460 83636 5470
rect 83580 5122 83636 5404
rect 83580 5070 83582 5122
rect 83634 5070 83636 5122
rect 83580 5058 83636 5070
rect 83468 5012 83524 5022
rect 83356 4900 83412 4910
rect 83356 4806 83412 4844
rect 83244 4286 83246 4338
rect 83298 4286 83300 4338
rect 83244 4274 83300 4286
rect 83356 4564 83412 4574
rect 83356 4338 83412 4508
rect 83356 4286 83358 4338
rect 83410 4286 83412 4338
rect 83356 4274 83412 4286
rect 83468 4340 83524 4956
rect 83692 4562 83748 7644
rect 83692 4510 83694 4562
rect 83746 4510 83748 4562
rect 83692 4498 83748 4510
rect 83804 4564 83860 9660
rect 83916 9650 83972 9660
rect 83916 7586 83972 7598
rect 83916 7534 83918 7586
rect 83970 7534 83972 7586
rect 83916 7364 83972 7534
rect 84028 7476 84084 12012
rect 84140 12002 84196 12012
rect 84812 12066 84868 20636
rect 86940 19236 86996 19246
rect 85932 18676 85988 18686
rect 84812 12014 84814 12066
rect 84866 12014 84868 12066
rect 84476 11172 84532 11182
rect 84476 11078 84532 11116
rect 84812 10724 84868 12014
rect 85372 13076 85428 13086
rect 85372 11508 85428 13020
rect 85932 12404 85988 18620
rect 84476 10668 84868 10724
rect 85260 11506 85428 11508
rect 85260 11454 85374 11506
rect 85426 11454 85428 11506
rect 85260 11452 85428 11454
rect 84252 8820 84308 8830
rect 84252 8258 84308 8764
rect 84252 8206 84254 8258
rect 84306 8206 84308 8258
rect 84252 8194 84308 8206
rect 84364 8034 84420 8046
rect 84364 7982 84366 8034
rect 84418 7982 84420 8034
rect 84364 7924 84420 7982
rect 84028 7410 84084 7420
rect 84252 7868 84420 7924
rect 83916 7298 83972 7308
rect 84028 7252 84084 7262
rect 83916 6580 83972 6590
rect 83916 5010 83972 6524
rect 84028 6018 84084 7196
rect 84140 6468 84196 6478
rect 84140 6374 84196 6412
rect 84028 5966 84030 6018
rect 84082 5966 84084 6018
rect 84028 5954 84084 5966
rect 83916 4958 83918 5010
rect 83970 4958 83972 5010
rect 83916 4946 83972 4958
rect 84140 5572 84196 5582
rect 84140 5012 84196 5516
rect 84252 5460 84308 7868
rect 84476 7812 84532 10668
rect 85260 10052 85316 11452
rect 85372 11442 85428 11452
rect 85484 12402 85988 12404
rect 85484 12350 85934 12402
rect 85986 12350 85988 12402
rect 85484 12348 85988 12350
rect 85484 10948 85540 12348
rect 85932 12272 85988 12348
rect 85260 9986 85316 9996
rect 85372 10892 85540 10948
rect 86380 10948 86436 10958
rect 84588 9940 84644 9950
rect 84588 9846 84644 9884
rect 84924 9716 84980 9726
rect 84812 8372 84868 8382
rect 84588 8258 84644 8270
rect 84588 8206 84590 8258
rect 84642 8206 84644 8258
rect 84588 8148 84644 8206
rect 84700 8148 84756 8158
rect 84588 8092 84700 8148
rect 84700 8082 84756 8092
rect 84252 5394 84308 5404
rect 84364 7756 84532 7812
rect 84252 5236 84308 5246
rect 84364 5236 84420 7756
rect 84812 7474 84868 8316
rect 84812 7422 84814 7474
rect 84866 7422 84868 7474
rect 84812 7410 84868 7422
rect 84476 6578 84532 6590
rect 84476 6526 84478 6578
rect 84530 6526 84532 6578
rect 84476 5348 84532 6526
rect 84476 5282 84532 5292
rect 84588 6468 84644 6478
rect 84252 5234 84420 5236
rect 84252 5182 84254 5234
rect 84306 5182 84420 5234
rect 84252 5180 84420 5182
rect 84252 5170 84308 5180
rect 84476 5124 84532 5134
rect 84364 5122 84532 5124
rect 84364 5070 84478 5122
rect 84530 5070 84532 5122
rect 84364 5068 84532 5070
rect 84364 5012 84420 5068
rect 84476 5058 84532 5068
rect 84140 4956 84420 5012
rect 84588 5012 84644 6412
rect 84028 4900 84084 4910
rect 84028 4806 84084 4844
rect 83804 4498 83860 4508
rect 84476 4788 84532 4798
rect 84476 4562 84532 4732
rect 84476 4510 84478 4562
rect 84530 4510 84532 4562
rect 84476 4498 84532 4510
rect 84588 4562 84644 4956
rect 84588 4510 84590 4562
rect 84642 4510 84644 4562
rect 84588 4498 84644 4510
rect 84700 5460 84756 5470
rect 84252 4452 84308 4462
rect 83580 4340 83636 4350
rect 83468 4338 83636 4340
rect 83468 4286 83582 4338
rect 83634 4286 83636 4338
rect 83468 4284 83636 4286
rect 83580 4274 83636 4284
rect 83804 4340 83860 4350
rect 82124 3502 82126 3554
rect 82178 3502 82180 3554
rect 82124 3490 82180 3502
rect 82796 3666 82852 3678
rect 82796 3614 82798 3666
rect 82850 3614 82852 3666
rect 82796 3388 82852 3614
rect 82012 1250 82068 1260
rect 82684 3332 82852 3388
rect 82684 800 82740 3332
rect 83804 2436 83860 4284
rect 84252 3554 84308 4396
rect 84700 4338 84756 5404
rect 84924 4900 84980 9660
rect 85148 9604 85204 9614
rect 85036 8596 85092 8606
rect 85036 8148 85092 8540
rect 85036 7586 85092 8092
rect 85036 7534 85038 7586
rect 85090 7534 85092 7586
rect 85036 7522 85092 7534
rect 84924 4834 84980 4844
rect 85036 5908 85092 5918
rect 84700 4286 84702 4338
rect 84754 4286 84756 4338
rect 84700 4274 84756 4286
rect 84812 4452 84868 4462
rect 84252 3502 84254 3554
rect 84306 3502 84308 3554
rect 84252 3490 84308 3502
rect 83804 2370 83860 2380
rect 84364 3444 84420 3454
rect 84364 800 84420 3388
rect 84812 1540 84868 4396
rect 85036 4450 85092 5852
rect 85148 5572 85204 9548
rect 85260 8146 85316 8158
rect 85260 8094 85262 8146
rect 85314 8094 85316 8146
rect 85260 8036 85316 8094
rect 85260 7970 85316 7980
rect 85260 6692 85316 6702
rect 85260 6598 85316 6636
rect 85148 5506 85204 5516
rect 85148 4564 85204 4574
rect 85148 4470 85204 4508
rect 85036 4398 85038 4450
rect 85090 4398 85092 4450
rect 85036 4386 85092 4398
rect 85372 4338 85428 10892
rect 86380 10834 86436 10892
rect 86380 10782 86382 10834
rect 86434 10782 86436 10834
rect 86380 10770 86436 10782
rect 86156 10610 86212 10622
rect 86156 10558 86158 10610
rect 86210 10558 86212 10610
rect 85596 10500 85652 10510
rect 85484 10498 85764 10500
rect 85484 10446 85598 10498
rect 85650 10446 85764 10498
rect 85484 10444 85764 10446
rect 85484 10388 85540 10444
rect 85596 10368 85652 10444
rect 85484 10322 85540 10332
rect 85484 9604 85540 9614
rect 85484 9602 85652 9604
rect 85484 9550 85486 9602
rect 85538 9550 85652 9602
rect 85484 9548 85652 9550
rect 85484 9538 85540 9548
rect 85484 8260 85540 8270
rect 85484 8166 85540 8204
rect 85484 6468 85540 6478
rect 85484 6374 85540 6412
rect 85596 6244 85652 9548
rect 85708 9156 85764 10444
rect 85708 9090 85764 9100
rect 85820 10052 85876 10062
rect 85820 9938 85876 9996
rect 85820 9886 85822 9938
rect 85874 9886 85876 9938
rect 85708 8930 85764 8942
rect 85708 8878 85710 8930
rect 85762 8878 85764 8930
rect 85708 8370 85764 8878
rect 85708 8318 85710 8370
rect 85762 8318 85764 8370
rect 85708 8306 85764 8318
rect 85820 8372 85876 9886
rect 86156 9492 86212 10558
rect 86492 10388 86548 10398
rect 86492 10386 86660 10388
rect 86492 10334 86494 10386
rect 86546 10334 86660 10386
rect 86492 10332 86660 10334
rect 86492 10322 86548 10332
rect 86492 9604 86548 9614
rect 86156 9426 86212 9436
rect 86380 9602 86548 9604
rect 86380 9550 86494 9602
rect 86546 9550 86548 9602
rect 86380 9548 86548 9550
rect 85820 8306 85876 8316
rect 86268 8372 86324 8382
rect 86268 8278 86324 8316
rect 85820 8146 85876 8158
rect 85820 8094 85822 8146
rect 85874 8094 85876 8146
rect 85820 6802 85876 8094
rect 86380 7588 86436 9548
rect 86492 9538 86548 9548
rect 86492 9044 86548 9054
rect 86492 8950 86548 8988
rect 85820 6750 85822 6802
rect 85874 6750 85876 6802
rect 85820 6738 85876 6750
rect 85932 7532 86436 7588
rect 86492 8148 86548 8158
rect 85820 6580 85876 6590
rect 85820 6486 85876 6524
rect 85596 6178 85652 6188
rect 85708 6466 85764 6478
rect 85708 6414 85710 6466
rect 85762 6414 85764 6466
rect 85708 6244 85764 6414
rect 85932 6244 85988 7532
rect 86492 7362 86548 8092
rect 86604 7812 86660 10332
rect 86940 10050 86996 19180
rect 86940 9998 86942 10050
rect 86994 9998 86996 10050
rect 86940 9938 86996 9998
rect 86940 9886 86942 9938
rect 86994 9886 86996 9938
rect 86940 9874 86996 9886
rect 87052 17780 87108 17790
rect 87052 10498 87108 17724
rect 88844 17668 88900 17678
rect 87836 15428 87892 15438
rect 87836 15148 87892 15372
rect 87836 15092 88004 15148
rect 87612 11282 87668 11294
rect 87612 11230 87614 11282
rect 87666 11230 87668 11282
rect 87612 10948 87668 11230
rect 87612 10882 87668 10892
rect 87052 10446 87054 10498
rect 87106 10446 87108 10498
rect 86940 8930 86996 8942
rect 86940 8878 86942 8930
rect 86994 8878 86996 8930
rect 86940 8372 86996 8878
rect 86828 8260 86884 8270
rect 86716 8148 86772 8158
rect 86716 8054 86772 8092
rect 86604 7756 86772 7812
rect 86492 7310 86494 7362
rect 86546 7310 86548 7362
rect 86492 7298 86548 7310
rect 85708 6188 85988 6244
rect 86380 6804 86436 6814
rect 85484 6020 85540 6030
rect 85484 5906 85540 5964
rect 85484 5854 85486 5906
rect 85538 5854 85540 5906
rect 85484 5842 85540 5854
rect 85596 5794 85652 5806
rect 85596 5742 85598 5794
rect 85650 5742 85652 5794
rect 85484 5236 85540 5246
rect 85484 5122 85540 5180
rect 85484 5070 85486 5122
rect 85538 5070 85540 5122
rect 85484 5058 85540 5070
rect 85596 4788 85652 5742
rect 85596 4722 85652 4732
rect 85372 4286 85374 4338
rect 85426 4286 85428 4338
rect 85372 4274 85428 4286
rect 85596 4340 85652 4350
rect 85596 4246 85652 4284
rect 85148 3444 85204 3482
rect 85148 3378 85204 3388
rect 84812 1474 84868 1484
rect 85708 1092 85764 6188
rect 86044 6020 86100 6030
rect 86044 5926 86100 5964
rect 85820 4900 85876 4910
rect 85820 4806 85876 4844
rect 86380 4450 86436 6748
rect 86716 6692 86772 7756
rect 86828 7474 86884 8204
rect 86940 8036 86996 8316
rect 86940 7970 86996 7980
rect 86828 7422 86830 7474
rect 86882 7422 86884 7474
rect 86828 7410 86884 7422
rect 86716 6626 86772 6636
rect 86828 6578 86884 6590
rect 86828 6526 86830 6578
rect 86882 6526 86884 6578
rect 86492 6468 86548 6478
rect 86492 6466 86660 6468
rect 86492 6414 86494 6466
rect 86546 6414 86660 6466
rect 86492 6412 86660 6414
rect 86492 6402 86548 6412
rect 86492 5796 86548 5806
rect 86492 5010 86548 5740
rect 86604 5460 86660 6412
rect 86828 6244 86884 6526
rect 87052 6580 87108 10446
rect 87612 10724 87668 10734
rect 87612 10498 87668 10668
rect 87612 10446 87614 10498
rect 87666 10446 87668 10498
rect 87612 10164 87668 10446
rect 87612 10098 87668 10108
rect 87164 10050 87220 10062
rect 87164 9998 87166 10050
rect 87218 9998 87220 10050
rect 87164 8428 87220 9998
rect 87500 10052 87556 10062
rect 87500 9602 87556 9996
rect 87612 9716 87668 9726
rect 87612 9622 87668 9660
rect 87724 9714 87780 9726
rect 87724 9662 87726 9714
rect 87778 9662 87780 9714
rect 87500 9550 87502 9602
rect 87554 9550 87556 9602
rect 87500 9492 87556 9550
rect 87500 9426 87556 9436
rect 87612 8930 87668 8942
rect 87612 8878 87614 8930
rect 87666 8878 87668 8930
rect 87164 8372 87444 8428
rect 87276 8260 87332 8270
rect 87276 8166 87332 8204
rect 87276 7364 87332 7374
rect 87052 6514 87108 6524
rect 87164 7362 87332 7364
rect 87164 7310 87278 7362
rect 87330 7310 87332 7362
rect 87164 7308 87332 7310
rect 86828 6178 86884 6188
rect 86604 5124 86660 5404
rect 86716 5124 86772 5134
rect 86604 5122 86772 5124
rect 86604 5070 86718 5122
rect 86770 5070 86772 5122
rect 86604 5068 86772 5070
rect 86716 5058 86772 5068
rect 87164 5122 87220 7308
rect 87276 7298 87332 7308
rect 87276 6804 87332 6814
rect 87276 6690 87332 6748
rect 87276 6638 87278 6690
rect 87330 6638 87332 6690
rect 87276 6626 87332 6638
rect 87388 5234 87444 8372
rect 87500 8258 87556 8270
rect 87500 8206 87502 8258
rect 87554 8206 87556 8258
rect 87500 8148 87556 8206
rect 87500 6914 87556 8092
rect 87500 6862 87502 6914
rect 87554 6862 87556 6914
rect 87500 6850 87556 6862
rect 87388 5182 87390 5234
rect 87442 5182 87444 5234
rect 87388 5170 87444 5182
rect 87500 6692 87556 6702
rect 87500 5234 87556 6636
rect 87500 5182 87502 5234
rect 87554 5182 87556 5234
rect 87500 5170 87556 5182
rect 87612 5234 87668 8878
rect 87724 7588 87780 9662
rect 87836 8148 87892 8158
rect 87836 8054 87892 8092
rect 87724 7522 87780 7532
rect 87724 7364 87780 7374
rect 87724 7270 87780 7308
rect 87724 6914 87780 6926
rect 87724 6862 87726 6914
rect 87778 6862 87780 6914
rect 87724 6802 87780 6862
rect 87724 6750 87726 6802
rect 87778 6750 87780 6802
rect 87724 6738 87780 6750
rect 87836 6468 87892 6478
rect 87836 6018 87892 6412
rect 87836 5966 87838 6018
rect 87890 5966 87892 6018
rect 87836 5954 87892 5966
rect 87612 5182 87614 5234
rect 87666 5182 87668 5234
rect 87164 5070 87166 5122
rect 87218 5070 87220 5122
rect 87164 5058 87220 5070
rect 86492 4958 86494 5010
rect 86546 4958 86548 5010
rect 86492 4946 86548 4958
rect 86604 4900 86660 4910
rect 86604 4806 86660 4844
rect 86380 4398 86382 4450
rect 86434 4398 86436 4450
rect 86380 4386 86436 4398
rect 86716 4450 86772 4462
rect 86716 4398 86718 4450
rect 86770 4398 86772 4450
rect 85708 1026 85764 1036
rect 86268 3666 86324 3678
rect 86268 3614 86270 3666
rect 86322 3614 86324 3666
rect 86268 980 86324 3614
rect 86716 3556 86772 4398
rect 87052 3556 87108 3566
rect 86716 3554 87108 3556
rect 86716 3502 87054 3554
rect 87106 3502 87108 3554
rect 86716 3500 87108 3502
rect 87052 3490 87108 3500
rect 86044 924 86324 980
rect 87612 980 87668 5182
rect 87948 5236 88004 15092
rect 88396 11394 88452 11406
rect 88396 11342 88398 11394
rect 88450 11342 88452 11394
rect 88396 11172 88452 11342
rect 88172 10610 88228 10622
rect 88172 10558 88174 10610
rect 88226 10558 88228 10610
rect 88172 10052 88228 10558
rect 88284 10500 88340 10510
rect 88284 10406 88340 10444
rect 88172 9986 88228 9996
rect 88284 10164 88340 10174
rect 88284 9828 88340 10108
rect 88060 9826 88340 9828
rect 88060 9774 88286 9826
rect 88338 9774 88340 9826
rect 88060 9772 88340 9774
rect 88060 9266 88116 9772
rect 88284 9762 88340 9772
rect 88060 9214 88062 9266
rect 88114 9214 88116 9266
rect 88060 9202 88116 9214
rect 88172 9156 88228 9166
rect 88172 6468 88228 9100
rect 88396 8932 88452 11116
rect 88508 10388 88564 10398
rect 88508 10386 88676 10388
rect 88508 10334 88510 10386
rect 88562 10334 88676 10386
rect 88508 10332 88676 10334
rect 88508 10322 88564 10332
rect 88508 8932 88564 8942
rect 88396 8876 88508 8932
rect 88508 8838 88564 8876
rect 88396 8036 88452 8046
rect 88172 6402 88228 6412
rect 88284 8034 88452 8036
rect 88284 7982 88398 8034
rect 88450 7982 88452 8034
rect 88284 7980 88452 7982
rect 88172 6020 88228 6030
rect 87948 5170 88004 5180
rect 88060 6018 88228 6020
rect 88060 5966 88174 6018
rect 88226 5966 88228 6018
rect 88060 5964 88228 5966
rect 86044 800 86100 924
rect 87612 914 87668 924
rect 87724 4226 87780 4238
rect 87724 4174 87726 4226
rect 87778 4174 87780 4226
rect 87724 800 87780 4174
rect 88060 3556 88116 5964
rect 88172 5954 88228 5964
rect 88172 5236 88228 5246
rect 88172 5142 88228 5180
rect 88284 4338 88340 7980
rect 88396 7970 88452 7980
rect 88508 7364 88564 7374
rect 88508 7270 88564 7308
rect 88396 6466 88452 6478
rect 88396 6414 88398 6466
rect 88450 6414 88452 6466
rect 88396 6356 88452 6414
rect 88396 6290 88452 6300
rect 88620 5124 88676 10332
rect 88732 8146 88788 8158
rect 88732 8094 88734 8146
rect 88786 8094 88788 8146
rect 88732 7364 88788 8094
rect 88732 7298 88788 7308
rect 88620 5058 88676 5068
rect 88732 6244 88788 6254
rect 88284 4286 88286 4338
rect 88338 4286 88340 4338
rect 88284 4274 88340 4286
rect 88396 4564 88452 4574
rect 88284 3668 88340 3678
rect 88396 3668 88452 4508
rect 88284 3666 88452 3668
rect 88284 3614 88286 3666
rect 88338 3614 88452 3666
rect 88284 3612 88452 3614
rect 88732 3666 88788 6188
rect 88844 4564 88900 17612
rect 89852 16100 89908 16110
rect 89852 15148 89908 16044
rect 89740 15092 89908 15148
rect 89516 12180 89572 12190
rect 89516 11508 89572 12124
rect 89292 11506 89572 11508
rect 89292 11454 89518 11506
rect 89570 11454 89572 11506
rect 89292 11452 89572 11454
rect 88956 11396 89012 11406
rect 88956 10164 89012 11340
rect 88956 10098 89012 10108
rect 89068 9716 89124 9726
rect 89068 9622 89124 9660
rect 89292 9268 89348 11452
rect 89516 11442 89572 11452
rect 89068 9212 89348 9268
rect 89516 10498 89572 10510
rect 89516 10446 89518 10498
rect 89570 10446 89572 10498
rect 89068 6468 89124 9212
rect 89404 9154 89460 9166
rect 89404 9102 89406 9154
rect 89458 9102 89460 9154
rect 89292 9042 89348 9054
rect 89292 8990 89294 9042
rect 89346 8990 89348 9042
rect 89292 8148 89348 8990
rect 89292 7476 89348 8092
rect 89404 8036 89460 9102
rect 89516 8260 89572 10446
rect 89628 9042 89684 9054
rect 89628 8990 89630 9042
rect 89682 8990 89684 9042
rect 89628 8596 89684 8990
rect 89628 8530 89684 8540
rect 89516 8194 89572 8204
rect 89404 7942 89460 7980
rect 89516 7476 89572 7486
rect 89740 7476 89796 15092
rect 91084 12290 91140 12302
rect 91084 12238 91086 12290
rect 91138 12238 91140 12290
rect 90412 12066 90468 12078
rect 90412 12014 90414 12066
rect 90466 12014 90468 12066
rect 90188 11956 90244 11966
rect 90188 9268 90244 11900
rect 90412 11732 90468 12014
rect 90412 11508 90468 11676
rect 90412 11442 90468 11452
rect 91084 11732 91140 12238
rect 91196 12180 91252 12190
rect 91196 12178 91476 12180
rect 91196 12126 91198 12178
rect 91250 12126 91476 12178
rect 91196 12124 91476 12126
rect 91196 12114 91252 12124
rect 91084 10612 91140 11676
rect 91084 10546 91140 10556
rect 91308 11954 91364 11966
rect 91308 11902 91310 11954
rect 91362 11902 91364 11954
rect 91308 9828 91364 11902
rect 91420 11508 91476 12124
rect 91532 11844 91588 25564
rect 96636 24332 96900 24342
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96636 24266 96900 24276
rect 96636 22764 96900 22774
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96636 22698 96900 22708
rect 96636 21196 96900 21206
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96636 21130 96900 21140
rect 98364 20188 98420 27244
rect 100716 24500 100772 24510
rect 99036 20916 99092 20926
rect 98364 20132 98644 20188
rect 96636 19628 96900 19638
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96636 19562 96900 19572
rect 94444 19124 94500 19134
rect 92204 17892 92260 17902
rect 91532 11778 91588 11788
rect 91756 13860 91812 13870
rect 91644 11508 91700 11518
rect 91420 11506 91700 11508
rect 91420 11454 91646 11506
rect 91698 11454 91700 11506
rect 91420 11452 91700 11454
rect 91644 11442 91700 11452
rect 91644 10500 91700 10510
rect 91644 10406 91700 10444
rect 91308 9772 91476 9828
rect 90188 9136 90244 9212
rect 91308 9602 91364 9614
rect 91308 9550 91310 9602
rect 91362 9550 91364 9602
rect 90300 8596 90356 8606
rect 90300 8370 90356 8540
rect 90300 8318 90302 8370
rect 90354 8318 90356 8370
rect 90300 8306 90356 8318
rect 90188 8260 90244 8270
rect 89292 7474 89572 7476
rect 89292 7422 89518 7474
rect 89570 7422 89572 7474
rect 89292 7420 89572 7422
rect 89516 7410 89572 7420
rect 89628 7420 89796 7476
rect 89852 8036 89908 8046
rect 89852 7474 89908 7980
rect 89852 7422 89854 7474
rect 89906 7422 89908 7474
rect 89628 7252 89684 7420
rect 89292 7196 89684 7252
rect 89292 6690 89348 7196
rect 89292 6638 89294 6690
rect 89346 6638 89348 6690
rect 89292 6626 89348 6638
rect 89068 6412 89348 6468
rect 88956 6356 89012 6366
rect 88956 5234 89012 6300
rect 89180 6244 89236 6254
rect 89180 6130 89236 6188
rect 89180 6078 89182 6130
rect 89234 6078 89236 6130
rect 89180 6066 89236 6078
rect 88956 5182 88958 5234
rect 89010 5182 89012 5234
rect 88956 5170 89012 5182
rect 89068 6020 89124 6030
rect 89068 5122 89124 5964
rect 89292 5908 89348 6412
rect 89068 5070 89070 5122
rect 89122 5070 89124 5122
rect 89068 5058 89124 5070
rect 89180 5852 89348 5908
rect 89628 5908 89684 7196
rect 89740 7252 89796 7262
rect 89740 6802 89796 7196
rect 89740 6750 89742 6802
rect 89794 6750 89796 6802
rect 89740 6738 89796 6750
rect 89852 6804 89908 7422
rect 90188 7252 90244 8204
rect 91084 8146 91140 8158
rect 91084 8094 91086 8146
rect 91138 8094 91140 8146
rect 90860 8036 90916 8046
rect 90860 7698 90916 7980
rect 90860 7646 90862 7698
rect 90914 7646 90916 7698
rect 90860 7634 90916 7646
rect 90748 7588 90804 7598
rect 90188 7186 90244 7196
rect 90412 7362 90468 7374
rect 90412 7310 90414 7362
rect 90466 7310 90468 7362
rect 89852 6738 89908 6748
rect 90076 6466 90132 6478
rect 90076 6414 90078 6466
rect 90130 6414 90132 6466
rect 90076 6244 90132 6414
rect 89740 5908 89796 5918
rect 89628 5906 89796 5908
rect 89628 5854 89742 5906
rect 89794 5854 89796 5906
rect 89628 5852 89796 5854
rect 88844 4498 88900 4508
rect 88732 3614 88734 3666
rect 88786 3614 88788 3666
rect 88284 3602 88340 3612
rect 88732 3602 88788 3614
rect 89180 4116 89236 5852
rect 89740 5842 89796 5852
rect 89964 5906 90020 5918
rect 89964 5854 89966 5906
rect 90018 5854 90020 5906
rect 89180 3666 89236 4060
rect 89180 3614 89182 3666
rect 89234 3614 89236 3666
rect 89180 3602 89236 3614
rect 89292 5348 89348 5358
rect 89292 4450 89348 5292
rect 89740 5012 89796 5022
rect 89740 4918 89796 4956
rect 89964 4900 90020 5854
rect 90076 5906 90132 6188
rect 90412 6018 90468 7310
rect 90524 6468 90580 6478
rect 90524 6374 90580 6412
rect 90412 5966 90414 6018
rect 90466 5966 90468 6018
rect 90412 5954 90468 5966
rect 90636 6244 90692 6254
rect 90076 5854 90078 5906
rect 90130 5854 90132 5906
rect 90076 5842 90132 5854
rect 90636 5460 90692 6188
rect 90748 6130 90804 7532
rect 90748 6078 90750 6130
rect 90802 6078 90804 6130
rect 90748 6066 90804 6078
rect 90972 6466 91028 6478
rect 90972 6414 90974 6466
rect 91026 6414 91028 6466
rect 90972 6020 91028 6414
rect 90972 5954 91028 5964
rect 90748 5908 90804 5918
rect 90748 5814 90804 5852
rect 90972 5796 91028 5806
rect 90972 5702 91028 5740
rect 91084 5572 91140 8094
rect 91308 8036 91364 9550
rect 91308 7970 91364 7980
rect 90300 5404 90692 5460
rect 89964 4834 90020 4844
rect 90188 4900 90244 4910
rect 90076 4564 90132 4574
rect 90076 4470 90132 4508
rect 90188 4562 90244 4844
rect 90188 4510 90190 4562
rect 90242 4510 90244 4562
rect 90188 4498 90244 4510
rect 89292 4398 89294 4450
rect 89346 4398 89348 4450
rect 88060 3490 88116 3500
rect 89292 1428 89348 4398
rect 89404 4340 89460 4350
rect 89404 4246 89460 4284
rect 90300 4338 90356 5404
rect 90412 5236 90468 5246
rect 90412 5010 90468 5180
rect 90636 5122 90692 5404
rect 90636 5070 90638 5122
rect 90690 5070 90692 5122
rect 90636 5058 90692 5070
rect 90748 5516 91140 5572
rect 91196 6914 91252 6926
rect 91196 6862 91198 6914
rect 91250 6862 91252 6914
rect 90412 4958 90414 5010
rect 90466 4958 90468 5010
rect 90412 4946 90468 4958
rect 90524 4900 90580 4910
rect 90748 4900 90804 5516
rect 91084 5124 91140 5134
rect 90972 5012 91028 5022
rect 90972 4918 91028 4956
rect 90524 4806 90580 4844
rect 90636 4844 90804 4900
rect 90636 4450 90692 4844
rect 91084 4562 91140 5068
rect 91084 4510 91086 4562
rect 91138 4510 91140 4562
rect 91084 4498 91140 4510
rect 90636 4398 90638 4450
rect 90690 4398 90692 4450
rect 90636 4386 90692 4398
rect 90300 4286 90302 4338
rect 90354 4286 90356 4338
rect 90300 4274 90356 4286
rect 91196 4338 91252 6862
rect 91308 5236 91364 5246
rect 91308 5142 91364 5180
rect 91420 5010 91476 9772
rect 91644 8372 91700 8382
rect 91644 8258 91700 8316
rect 91644 8206 91646 8258
rect 91698 8206 91700 8258
rect 91644 8194 91700 8206
rect 91756 7698 91812 13804
rect 92092 12292 92148 12302
rect 91868 8596 91924 8606
rect 91868 8370 91924 8540
rect 91868 8318 91870 8370
rect 91922 8318 91924 8370
rect 91868 8306 91924 8318
rect 91980 8148 92036 8158
rect 91980 8054 92036 8092
rect 92092 7924 92148 12236
rect 91756 7646 91758 7698
rect 91810 7646 91812 7698
rect 91756 6914 91812 7646
rect 91756 6862 91758 6914
rect 91810 6862 91812 6914
rect 91756 6850 91812 6862
rect 91980 7868 92148 7924
rect 91532 6692 91588 6702
rect 91532 5796 91588 6636
rect 91980 6690 92036 7868
rect 91980 6638 91982 6690
rect 92034 6638 92036 6690
rect 91868 6356 91924 6366
rect 91644 6020 91700 6030
rect 91644 5926 91700 5964
rect 91868 6018 91924 6300
rect 91868 5966 91870 6018
rect 91922 5966 91924 6018
rect 91868 5954 91924 5966
rect 91980 5908 92036 6638
rect 91980 5842 92036 5852
rect 92092 7362 92148 7374
rect 92092 7310 92094 7362
rect 92146 7310 92148 7362
rect 91532 5730 91588 5740
rect 91756 5796 91812 5806
rect 91756 5702 91812 5740
rect 91868 5572 91924 5582
rect 91644 5460 91700 5470
rect 91644 5234 91700 5404
rect 91644 5182 91646 5234
rect 91698 5182 91700 5234
rect 91644 5170 91700 5182
rect 91420 4958 91422 5010
rect 91474 4958 91476 5010
rect 91420 4946 91476 4958
rect 91308 4788 91364 4798
rect 91644 4788 91700 4798
rect 91364 4732 91644 4788
rect 91308 4722 91364 4732
rect 91644 4722 91700 4732
rect 91196 4286 91198 4338
rect 91250 4286 91252 4338
rect 91196 4274 91252 4286
rect 91756 4338 91812 4350
rect 91756 4286 91758 4338
rect 91810 4286 91812 4338
rect 90972 4228 91028 4238
rect 90972 4134 91028 4172
rect 91756 4116 91812 4286
rect 91756 4050 91812 4060
rect 89628 3556 89684 3566
rect 89628 3462 89684 3500
rect 89292 1362 89348 1372
rect 89404 3444 89460 3454
rect 89404 800 89460 3388
rect 90524 3444 90580 3482
rect 90524 3378 90580 3388
rect 91084 3444 91140 3454
rect 91084 800 91140 3388
rect 91868 2436 91924 5516
rect 92092 5348 92148 7310
rect 92092 5282 92148 5292
rect 92092 4900 92148 4910
rect 91980 4898 92148 4900
rect 91980 4846 92094 4898
rect 92146 4846 92148 4898
rect 91980 4844 92148 4846
rect 91980 4004 92036 4844
rect 92092 4834 92148 4844
rect 91980 3938 92036 3948
rect 92092 4450 92148 4462
rect 92092 4398 92094 4450
rect 92146 4398 92148 4450
rect 92092 3554 92148 4398
rect 92204 4228 92260 17836
rect 93436 15540 93492 15550
rect 92316 15428 92372 15438
rect 92316 6690 92372 15372
rect 93436 15148 93492 15484
rect 93324 15092 93492 15148
rect 92428 11396 92484 11406
rect 92428 10610 92484 11340
rect 92428 10558 92430 10610
rect 92482 10558 92484 10610
rect 92428 10546 92484 10558
rect 93212 9042 93268 9054
rect 93212 8990 93214 9042
rect 93266 8990 93268 9042
rect 92428 8930 92484 8942
rect 92428 8878 92430 8930
rect 92482 8878 92484 8930
rect 92428 8596 92484 8878
rect 93212 8932 93268 8990
rect 93212 8866 93268 8876
rect 92428 8530 92484 8540
rect 92988 8484 93044 8494
rect 92428 8372 92484 8382
rect 92428 8278 92484 8316
rect 92988 7700 93044 8428
rect 93100 8148 93156 8158
rect 93100 8036 93156 8092
rect 93100 8034 93268 8036
rect 93100 7982 93102 8034
rect 93154 7982 93268 8034
rect 93100 7980 93268 7982
rect 93100 7970 93156 7980
rect 93100 7700 93156 7710
rect 92988 7698 93156 7700
rect 92988 7646 93102 7698
rect 93154 7646 93156 7698
rect 92988 7644 93156 7646
rect 93100 7634 93156 7644
rect 92764 7364 92820 7374
rect 92316 6638 92318 6690
rect 92370 6638 92372 6690
rect 92316 5236 92372 6638
rect 92540 7362 92820 7364
rect 92540 7310 92766 7362
rect 92818 7310 92820 7362
rect 92540 7308 92820 7310
rect 92540 6244 92596 7308
rect 92764 7298 92820 7308
rect 93212 7252 93268 7980
rect 93212 7186 93268 7196
rect 93100 6692 93156 6702
rect 93324 6692 93380 15092
rect 93996 14756 94052 14766
rect 93660 12180 93716 12190
rect 92540 6178 92596 6188
rect 92652 6690 93380 6692
rect 92652 6638 93102 6690
rect 93154 6638 93380 6690
rect 92652 6636 93380 6638
rect 93548 11844 93604 11854
rect 93548 7700 93604 11788
rect 92540 6020 92596 6030
rect 92428 6018 92596 6020
rect 92428 5966 92542 6018
rect 92594 5966 92596 6018
rect 92428 5964 92596 5966
rect 92428 5460 92484 5964
rect 92540 5954 92596 5964
rect 92652 6018 92708 6636
rect 93100 6626 93156 6636
rect 93100 6356 93156 6366
rect 93100 6130 93156 6300
rect 93100 6078 93102 6130
rect 93154 6078 93156 6130
rect 93100 6066 93156 6078
rect 92652 5966 92654 6018
rect 92706 5966 92708 6018
rect 92652 5954 92708 5966
rect 92540 5684 92596 5694
rect 92540 5682 92708 5684
rect 92540 5630 92542 5682
rect 92594 5630 92708 5682
rect 92540 5628 92708 5630
rect 92540 5618 92596 5628
rect 92428 5404 92596 5460
rect 92316 5170 92372 5180
rect 92428 5010 92484 5022
rect 92428 4958 92430 5010
rect 92482 4958 92484 5010
rect 92428 4564 92484 4958
rect 92428 4498 92484 4508
rect 92540 4340 92596 5404
rect 92652 5348 92708 5628
rect 93324 5682 93380 5694
rect 93324 5630 93326 5682
rect 93378 5630 93380 5682
rect 92652 5292 92820 5348
rect 92764 4564 92820 5292
rect 93212 5012 93268 5022
rect 93212 4918 93268 4956
rect 92540 4274 92596 4284
rect 92652 4508 92820 4564
rect 93324 4564 93380 5630
rect 93548 5124 93604 7644
rect 93660 6130 93716 12124
rect 93772 11396 93828 11406
rect 93772 11302 93828 11340
rect 93996 9716 94052 14700
rect 94108 13972 94164 13982
rect 94108 10164 94164 13916
rect 94444 11788 94500 19068
rect 95564 19124 95620 19134
rect 95228 16324 95284 16334
rect 94780 16212 94836 16222
rect 94780 15148 94836 16156
rect 95228 15148 95284 16268
rect 94780 15092 94948 15148
rect 94444 11732 94612 11788
rect 94220 11396 94276 11406
rect 94276 11382 94388 11396
rect 94276 11340 94334 11382
rect 94220 11330 94276 11340
rect 94332 11330 94334 11340
rect 94386 11330 94388 11382
rect 94332 11318 94388 11330
rect 94108 10108 94500 10164
rect 93772 8484 93828 8494
rect 93772 8370 93828 8428
rect 93772 8318 93774 8370
rect 93826 8318 93828 8370
rect 93772 8306 93828 8318
rect 93996 7698 94052 9660
rect 94220 9156 94276 9166
rect 94220 8932 94276 9100
rect 94108 8930 94276 8932
rect 94108 8878 94222 8930
rect 94274 8878 94276 8930
rect 94108 8876 94276 8878
rect 94108 8484 94164 8876
rect 94220 8866 94276 8876
rect 94108 8418 94164 8428
rect 94220 8372 94276 8382
rect 94220 8278 94276 8316
rect 94444 7924 94500 10108
rect 94556 8148 94612 11732
rect 94668 9266 94724 9278
rect 94668 9214 94670 9266
rect 94722 9214 94724 9266
rect 94668 9156 94724 9214
rect 94780 9156 94836 9166
rect 94668 9154 94836 9156
rect 94668 9102 94782 9154
rect 94834 9102 94836 9154
rect 94668 9100 94836 9102
rect 94780 9090 94836 9100
rect 94892 8708 94948 15092
rect 95004 15092 95284 15148
rect 95004 10724 95060 15092
rect 95116 11282 95172 11294
rect 95116 11230 95118 11282
rect 95170 11230 95172 11282
rect 95116 10836 95172 11230
rect 95116 10780 95508 10836
rect 95004 10668 95284 10724
rect 95116 10500 95172 10510
rect 95004 9604 95060 9614
rect 95004 9510 95060 9548
rect 95004 9156 95060 9166
rect 95116 9156 95172 10444
rect 95004 9154 95172 9156
rect 95004 9102 95006 9154
rect 95058 9102 95118 9154
rect 95170 9102 95172 9154
rect 95004 9100 95172 9102
rect 95004 9090 95060 9100
rect 95116 9090 95172 9100
rect 94668 8652 94948 8708
rect 95228 8818 95284 10668
rect 95340 10276 95396 10286
rect 95340 9604 95396 10220
rect 95452 10050 95508 10780
rect 95452 9998 95454 10050
rect 95506 9998 95508 10050
rect 95452 9986 95508 9998
rect 95564 10052 95620 19068
rect 96636 18060 96900 18070
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96636 17994 96900 18004
rect 95564 9986 95620 9996
rect 95676 17444 95732 17454
rect 95564 9604 95620 9614
rect 95340 9602 95620 9604
rect 95340 9550 95566 9602
rect 95618 9550 95620 9602
rect 95340 9548 95620 9550
rect 95228 8766 95230 8818
rect 95282 8766 95284 8818
rect 94668 8260 94724 8652
rect 94780 8484 94836 8494
rect 94780 8390 94836 8428
rect 95228 8484 95284 8766
rect 94892 8260 94948 8270
rect 94668 8258 94948 8260
rect 94668 8206 94894 8258
rect 94946 8206 94948 8258
rect 94668 8204 94948 8206
rect 94556 8082 94612 8092
rect 94780 8036 94836 8046
rect 94444 7868 94612 7924
rect 93996 7646 93998 7698
rect 94050 7646 94052 7698
rect 93996 7588 94052 7646
rect 94444 7700 94500 7710
rect 94444 7606 94500 7644
rect 93996 7522 94052 7532
rect 93660 6078 93662 6130
rect 93714 6078 93716 6130
rect 93660 5460 93716 6078
rect 93660 5394 93716 5404
rect 93772 7476 93828 7486
rect 93772 6690 93828 7420
rect 93772 6638 93774 6690
rect 93826 6638 93828 6690
rect 93772 6132 93828 6638
rect 93772 5124 93828 6076
rect 94444 6466 94500 6478
rect 94444 6414 94446 6466
rect 94498 6414 94500 6466
rect 94444 5908 94500 6414
rect 94556 6356 94612 7868
rect 94780 7700 94836 7980
rect 94892 7924 94948 8204
rect 94892 7858 94948 7868
rect 95004 8148 95060 8158
rect 94892 7700 94948 7710
rect 94780 7698 94948 7700
rect 94780 7646 94894 7698
rect 94946 7646 94948 7698
rect 94780 7644 94948 7646
rect 94892 7634 94948 7644
rect 95004 7586 95060 8092
rect 95228 7812 95284 8428
rect 95340 8372 95396 8382
rect 95340 8278 95396 8316
rect 95452 8260 95508 9548
rect 95564 9538 95620 9548
rect 95676 9380 95732 17388
rect 97580 16884 97636 16894
rect 96636 16492 96900 16502
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96636 16426 96900 16436
rect 96348 15988 96404 15998
rect 96348 15148 96404 15932
rect 96124 15092 96404 15148
rect 97132 15876 97188 15886
rect 96012 11172 96068 11182
rect 96012 10498 96068 11116
rect 96012 10446 96014 10498
rect 96066 10446 96068 10498
rect 96012 10276 96068 10446
rect 96012 10210 96068 10220
rect 95788 9716 95844 9726
rect 95788 9714 96068 9716
rect 95788 9662 95790 9714
rect 95842 9662 96068 9714
rect 95788 9660 96068 9662
rect 95788 9650 95844 9660
rect 95676 9324 95844 9380
rect 95788 8372 95844 9324
rect 95788 8306 95844 8316
rect 95900 9042 95956 9054
rect 95900 8990 95902 9042
rect 95954 8990 95956 9042
rect 95452 8194 95508 8204
rect 95564 8258 95620 8270
rect 95564 8206 95566 8258
rect 95618 8206 95620 8258
rect 95564 8036 95620 8206
rect 95564 7970 95620 7980
rect 95676 8036 95732 8046
rect 95900 8036 95956 8990
rect 95676 8034 95956 8036
rect 95676 7982 95678 8034
rect 95730 7982 95956 8034
rect 95676 7980 95956 7982
rect 95676 7970 95732 7980
rect 95228 7746 95284 7756
rect 95340 7700 95396 7710
rect 95004 7534 95006 7586
rect 95058 7534 95060 7586
rect 95004 6804 95060 7534
rect 95228 7588 95284 7598
rect 95228 6916 95284 7532
rect 95340 7476 95396 7644
rect 95676 7588 95732 7598
rect 95452 7476 95508 7486
rect 95340 7474 95508 7476
rect 95340 7422 95454 7474
rect 95506 7422 95508 7474
rect 95340 7420 95508 7422
rect 95452 7410 95508 7420
rect 95228 6850 95284 6860
rect 95116 6804 95172 6814
rect 95004 6802 95172 6804
rect 95004 6750 95118 6802
rect 95170 6750 95172 6802
rect 95004 6748 95172 6750
rect 95116 6692 95172 6748
rect 95116 6626 95172 6636
rect 95676 6690 95732 7532
rect 96012 7140 96068 9660
rect 96124 7588 96180 15092
rect 96636 14924 96900 14934
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96636 14858 96900 14868
rect 96636 13356 96900 13366
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96636 13290 96900 13300
rect 96636 11788 96900 11798
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96636 11722 96900 11732
rect 97132 11732 97188 15820
rect 97132 11666 97188 11676
rect 97244 11508 97300 11518
rect 97580 11508 97636 16828
rect 98588 15148 98644 20132
rect 98588 15092 98756 15148
rect 98140 12066 98196 12078
rect 98140 12014 98142 12066
rect 98194 12014 98196 12066
rect 97132 11506 97636 11508
rect 97132 11454 97246 11506
rect 97298 11454 97636 11506
rect 97132 11452 97636 11454
rect 97692 11732 97748 11742
rect 96460 11396 96516 11406
rect 96460 10834 96516 11340
rect 96460 10782 96462 10834
rect 96514 10782 96516 10834
rect 96460 10770 96516 10782
rect 96636 10220 96900 10230
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96636 10154 96900 10164
rect 96572 9716 96628 9726
rect 96572 9622 96628 9660
rect 96908 9716 96964 9726
rect 97132 9716 97188 11452
rect 97244 11442 97300 11452
rect 97692 11172 97748 11676
rect 98140 11732 98196 12014
rect 98140 11396 98196 11676
rect 98140 11330 98196 11340
rect 98252 11172 98308 11182
rect 97692 11170 97860 11172
rect 97692 11118 97694 11170
rect 97746 11118 97860 11170
rect 97692 11116 97860 11118
rect 97692 11106 97748 11116
rect 97244 10500 97300 10510
rect 97244 10406 97300 10444
rect 97804 10500 97860 11116
rect 98252 11170 98532 11172
rect 98252 11118 98254 11170
rect 98306 11118 98532 11170
rect 98252 11116 98532 11118
rect 98252 11106 98308 11116
rect 97804 9828 97860 10444
rect 98252 10948 98308 10958
rect 98140 9828 98196 9838
rect 97804 9826 98196 9828
rect 97804 9774 98142 9826
rect 98194 9774 98196 9826
rect 97804 9772 98196 9774
rect 98140 9762 98196 9772
rect 96908 9714 97188 9716
rect 96908 9662 96910 9714
rect 96962 9662 97188 9714
rect 96908 9660 97188 9662
rect 97692 9714 97748 9726
rect 97692 9662 97694 9714
rect 97746 9662 97748 9714
rect 96908 9650 96964 9660
rect 96236 9268 96292 9278
rect 96236 9174 96292 9212
rect 96460 9154 96516 9166
rect 96460 9102 96462 9154
rect 96514 9102 96516 9154
rect 96348 8260 96404 8270
rect 96460 8260 96516 9102
rect 96572 8820 96628 8858
rect 96572 8754 96628 8764
rect 96636 8652 96900 8662
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96636 8586 96900 8596
rect 96684 8372 96740 8382
rect 96460 8204 96628 8260
rect 96348 8166 96404 8204
rect 96236 8036 96292 8046
rect 96236 7942 96292 7980
rect 96460 8034 96516 8046
rect 96460 7982 96462 8034
rect 96514 7982 96516 8034
rect 96460 7924 96516 7982
rect 96460 7858 96516 7868
rect 96572 7700 96628 8204
rect 96684 8146 96740 8316
rect 96684 8094 96686 8146
rect 96738 8094 96740 8146
rect 96684 8082 96740 8094
rect 96460 7644 96628 7700
rect 97020 7700 97076 9660
rect 97468 9604 97524 9614
rect 96124 7532 96404 7588
rect 96124 7364 96180 7374
rect 96124 7270 96180 7308
rect 96012 7084 96180 7140
rect 95676 6638 95678 6690
rect 95730 6638 95732 6690
rect 95676 6626 95732 6638
rect 95900 6692 95956 6730
rect 95900 6626 95956 6636
rect 95900 6466 95956 6478
rect 95900 6414 95902 6466
rect 95954 6414 95956 6466
rect 94556 6290 94612 6300
rect 95564 6356 95620 6366
rect 95004 6244 95060 6254
rect 95004 6132 95060 6188
rect 95004 6130 95172 6132
rect 95004 6078 95006 6130
rect 95058 6078 95172 6130
rect 95004 6076 95172 6078
rect 95004 6066 95060 6076
rect 94668 5908 94724 5918
rect 94444 5906 94724 5908
rect 94444 5854 94670 5906
rect 94722 5854 94724 5906
rect 94444 5852 94724 5854
rect 93996 5794 94052 5806
rect 93996 5742 93998 5794
rect 94050 5742 94052 5794
rect 93996 5682 94052 5742
rect 93996 5630 93998 5682
rect 94050 5630 94052 5682
rect 93996 5618 94052 5630
rect 93548 5068 93716 5124
rect 93660 5012 93716 5068
rect 93772 5058 93828 5068
rect 93660 4946 93716 4956
rect 94108 5012 94164 5022
rect 92204 4162 92260 4172
rect 92652 3780 92708 4508
rect 92988 4452 93044 4462
rect 92764 4340 92820 4350
rect 92764 4246 92820 4284
rect 92988 4338 93044 4396
rect 92988 4286 92990 4338
rect 93042 4286 93044 4338
rect 92988 4274 93044 4286
rect 92652 3714 92708 3724
rect 92092 3502 92094 3554
rect 92146 3502 92148 3554
rect 92092 3490 92148 3502
rect 92764 3556 92820 3566
rect 91868 2370 91924 2380
rect 92764 800 92820 3500
rect 92876 3444 92932 3482
rect 92876 3378 92932 3388
rect 93324 2772 93380 4508
rect 93548 4898 93604 4910
rect 93548 4846 93550 4898
rect 93602 4846 93604 4898
rect 93548 3556 93604 4846
rect 93772 4228 93828 4238
rect 93772 4134 93828 4172
rect 93772 3556 93828 3566
rect 93548 3554 93828 3556
rect 93548 3502 93774 3554
rect 93826 3502 93828 3554
rect 93548 3500 93828 3502
rect 93772 3490 93828 3500
rect 94108 3220 94164 4956
rect 94444 4898 94500 4910
rect 94444 4846 94446 4898
rect 94498 4846 94500 4898
rect 94444 4340 94500 4846
rect 94668 4900 94724 5852
rect 95004 5236 95060 5246
rect 95004 5010 95060 5180
rect 95004 4958 95006 5010
rect 95058 4958 95060 5010
rect 95004 4946 95060 4958
rect 94724 4844 94836 4900
rect 94668 4834 94724 4844
rect 94668 4340 94724 4350
rect 94444 4338 94724 4340
rect 94444 4286 94670 4338
rect 94722 4286 94724 4338
rect 94444 4284 94724 4286
rect 94668 4274 94724 4284
rect 94108 3154 94164 3164
rect 94444 3780 94500 3790
rect 93324 2706 93380 2716
rect 94444 800 94500 3724
rect 94780 3668 94836 4844
rect 95116 4564 95172 6076
rect 95564 6020 95620 6300
rect 95564 6018 95732 6020
rect 95564 5966 95566 6018
rect 95618 5966 95732 6018
rect 95564 5964 95732 5966
rect 95564 5954 95620 5964
rect 95340 4900 95396 4910
rect 95340 4806 95396 4844
rect 95116 4498 95172 4508
rect 95676 4452 95732 5964
rect 95788 5794 95844 5806
rect 95788 5742 95790 5794
rect 95842 5742 95844 5794
rect 95788 4564 95844 5742
rect 95900 5346 95956 6414
rect 96124 6130 96180 7084
rect 96236 6916 96292 6926
rect 96236 6692 96292 6860
rect 96236 6560 96292 6636
rect 96348 6244 96404 7532
rect 96460 6916 96516 7644
rect 97020 7634 97076 7644
rect 97132 9156 97188 9166
rect 96636 7084 96900 7094
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96636 7018 96900 7028
rect 96684 6916 96740 6926
rect 96460 6860 96684 6916
rect 96684 6802 96740 6860
rect 96684 6750 96686 6802
rect 96738 6750 96740 6802
rect 96684 6738 96740 6750
rect 96348 6188 97076 6244
rect 96124 6078 96126 6130
rect 96178 6078 96180 6130
rect 96124 6066 96180 6078
rect 96236 6020 96292 6030
rect 96236 5926 96292 5964
rect 96460 5908 96516 5918
rect 96348 5906 96516 5908
rect 96348 5854 96462 5906
rect 96514 5854 96516 5906
rect 96348 5852 96516 5854
rect 96012 5684 96068 5694
rect 96012 5590 96068 5628
rect 95900 5294 95902 5346
rect 95954 5294 95956 5346
rect 95900 5282 95956 5294
rect 96236 5348 96292 5358
rect 96348 5348 96404 5852
rect 96460 5842 96516 5852
rect 96636 5516 96900 5526
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96636 5450 96900 5460
rect 97020 5348 97076 6188
rect 96236 5346 96404 5348
rect 96236 5294 96238 5346
rect 96290 5294 96404 5346
rect 96236 5292 96404 5294
rect 96908 5292 97076 5348
rect 96236 5282 96292 5292
rect 96348 5124 96404 5134
rect 96124 5012 96180 5022
rect 96124 4918 96180 4956
rect 95788 4508 96292 4564
rect 95676 4396 95844 4452
rect 95340 4226 95396 4238
rect 95340 4174 95342 4226
rect 95394 4174 95396 4226
rect 95340 3780 95396 4174
rect 95340 3714 95396 3724
rect 94780 3602 94836 3612
rect 95788 3666 95844 4396
rect 95788 3614 95790 3666
rect 95842 3614 95844 3666
rect 95788 3602 95844 3614
rect 94668 3556 94724 3566
rect 94668 3462 94724 3500
rect 96124 3444 96180 3454
rect 96124 800 96180 3388
rect 96236 3332 96292 4508
rect 96348 4562 96404 5068
rect 96796 5012 96852 5022
rect 96348 4510 96350 4562
rect 96402 4510 96404 4562
rect 96348 4452 96404 4510
rect 96348 4386 96404 4396
rect 96460 4900 96516 4910
rect 96460 3554 96516 4844
rect 96796 4452 96852 4956
rect 96796 4386 96852 4396
rect 96908 5010 96964 5292
rect 96908 4958 96910 5010
rect 96962 4958 96964 5010
rect 96908 4116 96964 4958
rect 97132 5236 97188 9100
rect 97356 9156 97412 9166
rect 97356 9062 97412 9100
rect 97244 8818 97300 8830
rect 97244 8766 97246 8818
rect 97298 8766 97300 8818
rect 97244 8372 97300 8766
rect 97244 8306 97300 8316
rect 97244 8034 97300 8046
rect 97244 7982 97246 8034
rect 97298 7982 97300 8034
rect 97244 7700 97300 7982
rect 97244 7634 97300 7644
rect 97356 7924 97412 7934
rect 97356 7586 97412 7868
rect 97356 7534 97358 7586
rect 97410 7534 97412 7586
rect 97356 7522 97412 7534
rect 97468 7476 97524 9548
rect 97580 9602 97636 9614
rect 97580 9550 97582 9602
rect 97634 9550 97636 9602
rect 97580 9268 97636 9550
rect 97580 9202 97636 9212
rect 97692 9604 97748 9662
rect 97916 9604 97972 9614
rect 97692 8372 97748 9548
rect 97804 9602 97972 9604
rect 97804 9550 97918 9602
rect 97970 9550 97972 9602
rect 97804 9548 97972 9550
rect 97804 9380 97860 9548
rect 97916 9538 97972 9548
rect 98252 9380 98308 10892
rect 98364 9716 98420 9754
rect 98364 9650 98420 9660
rect 97804 9314 97860 9324
rect 97916 9324 98308 9380
rect 98364 9492 98420 9502
rect 97580 8316 97748 8372
rect 97580 7924 97636 8316
rect 97580 7858 97636 7868
rect 97804 8258 97860 8270
rect 97804 8206 97806 8258
rect 97858 8206 97860 8258
rect 97804 7924 97860 8206
rect 97804 7858 97860 7868
rect 97692 7812 97748 7822
rect 97692 7700 97748 7756
rect 97804 7700 97860 7710
rect 97692 7698 97860 7700
rect 97692 7646 97806 7698
rect 97858 7646 97860 7698
rect 97692 7644 97860 7646
rect 97804 7634 97860 7644
rect 97468 7420 97860 7476
rect 97244 7364 97300 7374
rect 97244 7270 97300 7308
rect 97580 7252 97636 7262
rect 97244 7028 97300 7038
rect 97244 6578 97300 6972
rect 97244 6526 97246 6578
rect 97298 6526 97300 6578
rect 97244 6514 97300 6526
rect 97356 6802 97412 6814
rect 97356 6750 97358 6802
rect 97410 6750 97412 6802
rect 97356 6020 97412 6750
rect 97468 6692 97524 6702
rect 97468 6598 97524 6636
rect 97356 5908 97412 5964
rect 97468 5908 97524 5918
rect 97356 5906 97524 5908
rect 97356 5854 97470 5906
rect 97522 5854 97524 5906
rect 97356 5852 97524 5854
rect 97468 5842 97524 5852
rect 97132 5122 97188 5180
rect 97132 5070 97134 5122
rect 97186 5070 97188 5122
rect 97020 4900 97076 4910
rect 97020 4564 97076 4844
rect 97132 4788 97188 5070
rect 97356 5682 97412 5694
rect 97356 5630 97358 5682
rect 97410 5630 97412 5682
rect 97356 5012 97412 5630
rect 97468 5012 97524 5022
rect 97356 5010 97524 5012
rect 97356 4958 97470 5010
rect 97522 4958 97524 5010
rect 97356 4956 97524 4958
rect 97468 4946 97524 4956
rect 97580 4898 97636 7196
rect 97692 6804 97748 6814
rect 97692 6690 97748 6748
rect 97692 6638 97694 6690
rect 97746 6638 97748 6690
rect 97692 6626 97748 6638
rect 97804 5236 97860 7420
rect 97580 4846 97582 4898
rect 97634 4846 97636 4898
rect 97580 4834 97636 4846
rect 97692 5234 97860 5236
rect 97692 5182 97806 5234
rect 97858 5182 97860 5234
rect 97692 5180 97860 5182
rect 97916 5236 97972 9324
rect 98252 9156 98308 9166
rect 98252 8820 98308 9100
rect 98364 9042 98420 9436
rect 98364 8990 98366 9042
rect 98418 8990 98420 9042
rect 98364 8978 98420 8990
rect 98252 8764 98420 8820
rect 98028 8146 98084 8158
rect 98028 8094 98030 8146
rect 98082 8094 98084 8146
rect 98028 7700 98084 8094
rect 98028 7634 98084 7644
rect 98140 8146 98196 8158
rect 98140 8094 98142 8146
rect 98194 8094 98196 8146
rect 98140 7588 98196 8094
rect 98140 7252 98196 7532
rect 98140 5906 98196 7196
rect 98252 7924 98308 7934
rect 98252 7140 98308 7868
rect 98364 7698 98420 8764
rect 98364 7646 98366 7698
rect 98418 7646 98420 7698
rect 98364 7634 98420 7646
rect 98252 7074 98308 7084
rect 98140 5854 98142 5906
rect 98194 5854 98196 5906
rect 98140 5842 98196 5854
rect 98252 6466 98308 6478
rect 98252 6414 98254 6466
rect 98306 6414 98308 6466
rect 98028 5236 98084 5246
rect 97916 5234 98084 5236
rect 97916 5182 98030 5234
rect 98082 5182 98084 5234
rect 97916 5180 98084 5182
rect 97132 4732 97524 4788
rect 97020 4498 97076 4508
rect 97356 4452 97412 4462
rect 97356 4358 97412 4396
rect 97468 4450 97524 4732
rect 97468 4398 97470 4450
rect 97522 4398 97524 4450
rect 97468 4386 97524 4398
rect 96908 4050 96964 4060
rect 96636 3948 96900 3958
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96636 3882 96900 3892
rect 96460 3502 96462 3554
rect 96514 3502 96516 3554
rect 96460 3490 96516 3502
rect 97244 3444 97300 3482
rect 97244 3378 97300 3388
rect 96236 3266 96292 3276
rect 97692 1652 97748 5180
rect 97804 5170 97860 5180
rect 98028 5170 98084 5180
rect 98252 4338 98308 6414
rect 98476 5124 98532 11116
rect 98700 10164 98756 15092
rect 98812 12178 98868 12190
rect 98812 12126 98814 12178
rect 98866 12126 98868 12178
rect 98812 11732 98868 12126
rect 98812 11666 98868 11676
rect 99036 10948 99092 20860
rect 100604 14532 100660 14542
rect 100492 13972 100548 13982
rect 100380 12740 100436 12750
rect 100156 12684 100380 12740
rect 99484 12068 99540 12078
rect 99260 12066 99540 12068
rect 99260 12014 99486 12066
rect 99538 12014 99540 12066
rect 99260 12012 99540 12014
rect 99260 11506 99316 12012
rect 99484 12002 99540 12012
rect 100156 11732 100212 12684
rect 100380 12608 100436 12684
rect 99260 11454 99262 11506
rect 99314 11454 99316 11506
rect 99260 11442 99316 11454
rect 99820 11618 99876 11630
rect 99820 11566 99822 11618
rect 99874 11566 99876 11618
rect 99372 11284 99428 11294
rect 99260 11282 99428 11284
rect 99260 11230 99374 11282
rect 99426 11230 99428 11282
rect 99260 11228 99428 11230
rect 99148 11172 99204 11182
rect 99148 11078 99204 11116
rect 99036 10882 99092 10892
rect 98588 8258 98644 8270
rect 98588 8206 98590 8258
rect 98642 8206 98644 8258
rect 98588 7476 98644 8206
rect 98700 7588 98756 10108
rect 98812 9826 98868 9838
rect 98812 9774 98814 9826
rect 98866 9774 98868 9826
rect 98812 9716 98868 9774
rect 98812 9042 98868 9660
rect 99148 9828 99204 9838
rect 99148 9380 99204 9772
rect 99148 9314 99204 9324
rect 98812 8990 98814 9042
rect 98866 8990 98868 9042
rect 98812 8482 98868 8990
rect 98812 8430 98814 8482
rect 98866 8430 98868 8482
rect 98812 8418 98868 8430
rect 98924 8930 98980 8942
rect 98924 8878 98926 8930
rect 98978 8878 98980 8930
rect 98700 7532 98868 7588
rect 98588 6804 98644 7420
rect 98700 7364 98756 7374
rect 98700 7270 98756 7308
rect 98588 6738 98644 6748
rect 98588 6580 98644 6590
rect 98812 6580 98868 7532
rect 98588 6578 98868 6580
rect 98588 6526 98590 6578
rect 98642 6526 98868 6578
rect 98588 6524 98868 6526
rect 98588 6514 98644 6524
rect 98924 6132 98980 8878
rect 99260 8484 99316 11228
rect 99372 11218 99428 11228
rect 99372 10500 99428 10510
rect 99372 10498 99764 10500
rect 99372 10446 99374 10498
rect 99426 10446 99764 10498
rect 99372 10444 99764 10446
rect 99372 10434 99428 10444
rect 99372 9604 99428 9614
rect 99372 9510 99428 9548
rect 99484 9604 99540 9614
rect 99484 9602 99652 9604
rect 99484 9550 99486 9602
rect 99538 9550 99652 9602
rect 99484 9548 99652 9550
rect 99484 9538 99540 9548
rect 99484 9156 99540 9166
rect 99484 9062 99540 9100
rect 99260 8428 99428 8484
rect 99148 8260 99204 8270
rect 99148 8166 99204 8204
rect 99260 8148 99316 8158
rect 99148 7364 99204 7374
rect 99148 7270 99204 7308
rect 99260 6916 99316 8092
rect 99036 6580 99092 6590
rect 99036 6486 99092 6524
rect 98924 6076 99092 6132
rect 98924 5908 98980 5918
rect 98924 5236 98980 5852
rect 98588 5124 98644 5134
rect 98476 5122 98644 5124
rect 98476 5070 98590 5122
rect 98642 5070 98644 5122
rect 98476 5068 98644 5070
rect 98476 4676 98532 5068
rect 98588 5058 98644 5068
rect 98812 5124 98868 5134
rect 98812 5010 98868 5068
rect 98924 5122 98980 5180
rect 98924 5070 98926 5122
rect 98978 5070 98980 5122
rect 98924 5058 98980 5070
rect 98812 4958 98814 5010
rect 98866 4958 98868 5010
rect 98812 4900 98868 4958
rect 99036 5012 99092 6076
rect 99260 6130 99316 6860
rect 99260 6078 99262 6130
rect 99314 6078 99316 6130
rect 99260 6066 99316 6078
rect 99260 5012 99316 5022
rect 99036 5010 99316 5012
rect 99036 4958 99262 5010
rect 99314 4958 99316 5010
rect 99036 4956 99316 4958
rect 99260 4946 99316 4956
rect 98812 4834 98868 4844
rect 99372 4898 99428 8428
rect 99484 8260 99540 8270
rect 99596 8260 99652 9548
rect 99708 9268 99764 10444
rect 99820 9828 99876 11566
rect 99932 11284 99988 11294
rect 99932 11190 99988 11228
rect 100044 11060 100100 11070
rect 99820 9772 99988 9828
rect 99820 9604 99876 9614
rect 99820 9510 99876 9548
rect 99820 9268 99876 9278
rect 99708 9266 99876 9268
rect 99708 9214 99822 9266
rect 99874 9214 99876 9266
rect 99708 9212 99876 9214
rect 99820 9202 99876 9212
rect 99932 9156 99988 9772
rect 99932 9090 99988 9100
rect 99708 9042 99764 9054
rect 99708 8990 99710 9042
rect 99762 8990 99764 9042
rect 99708 8820 99764 8990
rect 99708 8754 99764 8764
rect 100044 8596 100100 11004
rect 100156 10612 100212 11676
rect 100156 10518 100212 10556
rect 100268 11956 100324 11966
rect 100268 9940 100324 11900
rect 100380 11170 100436 11182
rect 100380 11118 100382 11170
rect 100434 11118 100436 11170
rect 100380 10948 100436 11118
rect 100380 10882 100436 10892
rect 100492 10164 100548 13916
rect 100604 11618 100660 14476
rect 100604 11566 100606 11618
rect 100658 11566 100660 11618
rect 100604 10834 100660 11566
rect 100716 11172 100772 24444
rect 100716 11106 100772 11116
rect 101052 11396 101108 115388
rect 102396 30324 102452 30334
rect 102060 21476 102116 21486
rect 101276 19012 101332 19022
rect 101164 12962 101220 12974
rect 101164 12910 101166 12962
rect 101218 12910 101220 12962
rect 101164 12740 101220 12910
rect 101164 12674 101220 12684
rect 101052 10836 101108 11340
rect 101164 11172 101220 11182
rect 101164 11078 101220 11116
rect 100604 10782 100606 10834
rect 100658 10782 100660 10834
rect 100604 10770 100660 10782
rect 100828 10834 101108 10836
rect 100828 10782 101054 10834
rect 101106 10782 101108 10834
rect 100828 10780 101108 10782
rect 100492 10108 100772 10164
rect 100268 9938 100548 9940
rect 100268 9886 100270 9938
rect 100322 9886 100548 9938
rect 100268 9884 100548 9886
rect 100268 9828 100324 9884
rect 100268 9762 100324 9772
rect 100380 9604 100436 9614
rect 100156 9044 100212 9054
rect 100156 9042 100324 9044
rect 100156 8990 100158 9042
rect 100210 8990 100324 9042
rect 100156 8988 100324 8990
rect 100156 8978 100212 8988
rect 99932 8540 100100 8596
rect 99484 8258 99652 8260
rect 99484 8206 99486 8258
rect 99538 8206 99652 8258
rect 99484 8204 99652 8206
rect 99708 8260 99764 8270
rect 99484 8194 99540 8204
rect 99708 8146 99764 8204
rect 99708 8094 99710 8146
rect 99762 8094 99764 8146
rect 99708 8082 99764 8094
rect 99820 8148 99876 8158
rect 99820 8054 99876 8092
rect 99932 7924 99988 8540
rect 99820 7868 99988 7924
rect 100044 8370 100100 8382
rect 100044 8318 100046 8370
rect 100098 8318 100100 8370
rect 99596 7812 99652 7822
rect 99484 6692 99540 6702
rect 99484 6598 99540 6636
rect 99596 5234 99652 7756
rect 99708 7700 99764 7710
rect 99708 7606 99764 7644
rect 99820 6244 99876 7868
rect 100044 7698 100100 8318
rect 100156 8372 100212 8382
rect 100156 8278 100212 8316
rect 100044 7646 100046 7698
rect 100098 7646 100100 7698
rect 100044 7634 100100 7646
rect 100156 8036 100212 8046
rect 100156 6916 100212 7980
rect 99932 6692 99988 6702
rect 99932 6598 99988 6636
rect 99596 5182 99598 5234
rect 99650 5182 99652 5234
rect 99596 5170 99652 5182
rect 99708 6188 99876 6244
rect 99372 4846 99374 4898
rect 99426 4846 99428 4898
rect 99372 4834 99428 4846
rect 98476 4610 98532 4620
rect 99708 4452 99764 6188
rect 99820 6020 99876 6030
rect 99820 6018 99988 6020
rect 99820 5966 99822 6018
rect 99874 5966 99988 6018
rect 99820 5964 99988 5966
rect 99820 5954 99876 5964
rect 99820 5236 99876 5246
rect 99820 5142 99876 5180
rect 99820 4452 99876 4462
rect 99708 4450 99876 4452
rect 99708 4398 99822 4450
rect 99874 4398 99876 4450
rect 99708 4396 99876 4398
rect 99820 4386 99876 4396
rect 98252 4286 98254 4338
rect 98306 4286 98308 4338
rect 98252 4274 98308 4286
rect 97692 1586 97748 1596
rect 97804 4228 97860 4238
rect 97804 800 97860 4172
rect 98700 4228 98756 4238
rect 98700 4134 98756 4172
rect 98924 4116 98980 4126
rect 98924 3666 98980 4060
rect 98924 3614 98926 3666
rect 98978 3614 98980 3666
rect 98924 3602 98980 3614
rect 98476 3556 98532 3566
rect 98476 3462 98532 3500
rect 99932 3554 99988 5964
rect 100156 6018 100212 6860
rect 100156 5966 100158 6018
rect 100210 5966 100212 6018
rect 100156 5954 100212 5966
rect 100268 5684 100324 8988
rect 100380 8482 100436 9548
rect 100492 9266 100548 9884
rect 100492 9214 100494 9266
rect 100546 9214 100548 9266
rect 100492 9202 100548 9214
rect 100604 9156 100660 9166
rect 100380 8430 100382 8482
rect 100434 8430 100436 8482
rect 100380 8418 100436 8430
rect 100492 8708 100548 8718
rect 100492 7812 100548 8652
rect 100604 8260 100660 9100
rect 100604 8194 100660 8204
rect 100492 7746 100548 7756
rect 100492 7476 100548 7486
rect 100492 7382 100548 7420
rect 100380 7364 100436 7374
rect 100380 6468 100436 7308
rect 100380 6466 100548 6468
rect 100380 6414 100382 6466
rect 100434 6414 100548 6466
rect 100380 6412 100548 6414
rect 100380 6402 100436 6412
rect 100156 5628 100324 5684
rect 100156 4562 100212 5628
rect 100268 5460 100324 5470
rect 100268 5234 100324 5404
rect 100268 5182 100270 5234
rect 100322 5182 100324 5234
rect 100268 5170 100324 5182
rect 100380 5012 100436 5022
rect 100156 4510 100158 4562
rect 100210 4510 100212 4562
rect 100156 4498 100212 4510
rect 100268 4676 100324 4686
rect 100268 4562 100324 4620
rect 100268 4510 100270 4562
rect 100322 4510 100324 4562
rect 100268 4498 100324 4510
rect 100380 4562 100436 4956
rect 100380 4510 100382 4562
rect 100434 4510 100436 4562
rect 100380 4498 100436 4510
rect 99932 3502 99934 3554
rect 99986 3502 99988 3554
rect 99932 3490 99988 3502
rect 100044 4338 100100 4350
rect 100044 4286 100046 4338
rect 100098 4286 100100 4338
rect 99484 3444 99540 3454
rect 98140 3332 98196 3342
rect 98140 3238 98196 3276
rect 98588 1652 98644 1662
rect 5936 0 6048 800
rect 6496 0 6608 800
rect 7056 0 7168 800
rect 7616 0 7728 800
rect 8176 0 8288 800
rect 8736 0 8848 800
rect 9296 0 9408 800
rect 9856 0 9968 800
rect 10416 0 10528 800
rect 10976 0 11088 800
rect 11536 0 11648 800
rect 12096 0 12208 800
rect 12656 0 12768 800
rect 13216 0 13328 800
rect 13776 0 13888 800
rect 14336 0 14448 800
rect 14896 0 15008 800
rect 15456 0 15568 800
rect 16016 0 16128 800
rect 16576 0 16688 800
rect 17136 0 17248 800
rect 17696 0 17808 800
rect 18256 0 18368 800
rect 18816 0 18928 800
rect 19376 0 19488 800
rect 19936 0 20048 800
rect 20496 0 20608 800
rect 21056 0 21168 800
rect 21616 0 21728 800
rect 22176 0 22288 800
rect 22736 0 22848 800
rect 23296 0 23408 800
rect 23856 0 23968 800
rect 24416 0 24528 800
rect 24976 0 25088 800
rect 25536 0 25648 800
rect 26096 0 26208 800
rect 26656 0 26768 800
rect 27216 0 27328 800
rect 27776 0 27888 800
rect 28336 0 28448 800
rect 28896 0 29008 800
rect 29456 0 29568 800
rect 30016 0 30128 800
rect 30576 0 30688 800
rect 31136 0 31248 800
rect 31696 0 31808 800
rect 32256 0 32368 800
rect 32816 0 32928 800
rect 33376 0 33488 800
rect 33936 0 34048 800
rect 34496 0 34608 800
rect 35056 0 35168 800
rect 35616 0 35728 800
rect 36176 0 36288 800
rect 36736 0 36848 800
rect 37296 0 37408 800
rect 37856 0 37968 800
rect 38416 0 38528 800
rect 38976 0 39088 800
rect 39536 0 39648 800
rect 40096 0 40208 800
rect 40656 0 40768 800
rect 41216 0 41328 800
rect 41776 0 41888 800
rect 42336 0 42448 800
rect 42896 0 43008 800
rect 43456 0 43568 800
rect 44016 0 44128 800
rect 44576 0 44688 800
rect 45136 0 45248 800
rect 45696 0 45808 800
rect 46256 0 46368 800
rect 46816 0 46928 800
rect 47376 0 47488 800
rect 47936 0 48048 800
rect 48496 0 48608 800
rect 49056 0 49168 800
rect 49616 0 49728 800
rect 50176 0 50288 800
rect 50736 0 50848 800
rect 51296 0 51408 800
rect 51856 0 51968 800
rect 52416 0 52528 800
rect 52976 0 53088 800
rect 53536 0 53648 800
rect 54096 0 54208 800
rect 54656 0 54768 800
rect 55216 0 55328 800
rect 55776 0 55888 800
rect 56336 0 56448 800
rect 56896 0 57008 800
rect 57456 0 57568 800
rect 58016 0 58128 800
rect 58576 0 58688 800
rect 59136 0 59248 800
rect 59696 0 59808 800
rect 60256 0 60368 800
rect 60816 0 60928 800
rect 61376 0 61488 800
rect 61936 0 62048 800
rect 62496 0 62608 800
rect 63056 0 63168 800
rect 63616 0 63728 800
rect 64176 0 64288 800
rect 64736 0 64848 800
rect 65296 0 65408 800
rect 65856 0 65968 800
rect 66416 0 66528 800
rect 66976 0 67088 800
rect 67536 0 67648 800
rect 68096 0 68208 800
rect 68656 0 68768 800
rect 69216 0 69328 800
rect 69776 0 69888 800
rect 70336 0 70448 800
rect 70896 0 71008 800
rect 71456 0 71568 800
rect 72016 0 72128 800
rect 72576 0 72688 800
rect 73136 0 73248 800
rect 73696 0 73808 800
rect 74256 0 74368 800
rect 74816 0 74928 800
rect 75376 0 75488 800
rect 75936 0 76048 800
rect 76496 0 76608 800
rect 77056 0 77168 800
rect 77616 0 77728 800
rect 78176 0 78288 800
rect 78736 0 78848 800
rect 79296 0 79408 800
rect 79856 0 79968 800
rect 80416 0 80528 800
rect 80976 0 81088 800
rect 81536 0 81648 800
rect 82096 0 82208 800
rect 82656 0 82768 800
rect 83216 0 83328 800
rect 83776 0 83888 800
rect 84336 0 84448 800
rect 84896 0 85008 800
rect 85456 0 85568 800
rect 86016 0 86128 800
rect 86576 0 86688 800
rect 87136 0 87248 800
rect 87696 0 87808 800
rect 88256 0 88368 800
rect 88816 0 88928 800
rect 89376 0 89488 800
rect 89936 0 90048 800
rect 90496 0 90608 800
rect 91056 0 91168 800
rect 91616 0 91728 800
rect 92176 0 92288 800
rect 92736 0 92848 800
rect 93296 0 93408 800
rect 93856 0 93968 800
rect 94416 0 94528 800
rect 94976 0 95088 800
rect 95536 0 95648 800
rect 96096 0 96208 800
rect 96656 0 96768 800
rect 97216 0 97328 800
rect 97776 0 97888 800
rect 98336 0 98448 800
rect 98588 756 98644 1596
rect 99484 800 99540 3388
rect 100044 3332 100100 4286
rect 100044 3266 100100 3276
rect 100492 1428 100548 6412
rect 100716 6130 100772 10108
rect 100828 8036 100884 10780
rect 101052 10770 101108 10780
rect 101276 10388 101332 18956
rect 102060 15148 102116 21420
rect 101836 15092 102116 15148
rect 101836 12628 101892 15092
rect 101948 12852 102004 12862
rect 101948 12850 102228 12852
rect 101948 12798 101950 12850
rect 102002 12798 102228 12850
rect 101948 12796 102228 12798
rect 101948 12786 102004 12796
rect 101836 12572 102004 12628
rect 101612 12066 101668 12078
rect 101612 12014 101614 12066
rect 101666 12014 101668 12066
rect 101612 11396 101668 12014
rect 101164 10386 101332 10388
rect 101164 10334 101278 10386
rect 101330 10334 101332 10386
rect 101164 10332 101332 10334
rect 101052 9716 101108 9726
rect 100940 9714 101108 9716
rect 100940 9662 101054 9714
rect 101106 9662 101108 9714
rect 100940 9660 101108 9662
rect 100940 9604 100996 9660
rect 101052 9650 101108 9660
rect 100940 9268 100996 9548
rect 100940 9174 100996 9212
rect 100828 7970 100884 7980
rect 100940 7700 100996 7710
rect 100940 7606 100996 7644
rect 101052 7476 101108 7486
rect 101052 6690 101108 7420
rect 101052 6638 101054 6690
rect 101106 6638 101108 6690
rect 101052 6626 101108 6638
rect 100716 6078 100718 6130
rect 100770 6078 100772 6130
rect 100716 5684 100772 6078
rect 100716 5618 100772 5628
rect 101164 6020 101220 10332
rect 101276 10322 101332 10332
rect 101388 11340 101668 11396
rect 101724 11396 101780 11406
rect 101388 10164 101444 11340
rect 101724 11284 101780 11340
rect 101612 11228 101780 11284
rect 101500 11170 101556 11182
rect 101500 11118 101502 11170
rect 101554 11118 101556 11170
rect 101500 11060 101556 11118
rect 101500 10994 101556 11004
rect 101276 10108 101444 10164
rect 101612 10834 101668 11228
rect 101948 11170 102004 12572
rect 101948 11118 101950 11170
rect 102002 11118 102004 11170
rect 101948 10836 102004 11118
rect 101612 10782 101614 10834
rect 101666 10782 101668 10834
rect 101276 9604 101332 10108
rect 101500 9604 101556 9614
rect 101276 9538 101332 9548
rect 101388 9602 101556 9604
rect 101388 9550 101502 9602
rect 101554 9550 101556 9602
rect 101388 9548 101556 9550
rect 101388 9044 101444 9548
rect 101500 9538 101556 9548
rect 101388 8978 101444 8988
rect 101500 8930 101556 8942
rect 101500 8878 101502 8930
rect 101554 8878 101556 8930
rect 101052 5236 101108 5246
rect 101052 5142 101108 5180
rect 101052 4564 101108 4574
rect 101164 4564 101220 5964
rect 101276 8484 101332 8494
rect 101276 5906 101332 8428
rect 101388 8260 101444 8270
rect 101388 8166 101444 8204
rect 101500 7924 101556 8878
rect 101612 8708 101668 10782
rect 101612 8642 101668 8652
rect 101724 10780 102004 10836
rect 101612 8148 101668 8158
rect 101612 8054 101668 8092
rect 101500 7858 101556 7868
rect 101500 7700 101556 7710
rect 101500 6802 101556 7644
rect 101500 6750 101502 6802
rect 101554 6750 101556 6802
rect 101500 6738 101556 6750
rect 101724 6580 101780 10780
rect 102172 10724 102228 12796
rect 101836 10668 102228 10724
rect 101836 8370 101892 10668
rect 101948 10498 102004 10510
rect 102396 10500 102452 30268
rect 104412 25508 104468 25518
rect 104300 21364 104356 21374
rect 104076 13074 104132 13086
rect 104076 13022 104078 13074
rect 104130 13022 104132 13074
rect 104076 11956 104132 13022
rect 104076 11890 104132 11900
rect 104300 11508 104356 21308
rect 104300 11442 104356 11452
rect 103404 11394 103460 11406
rect 103404 11342 103406 11394
rect 103458 11342 103460 11394
rect 101948 10446 101950 10498
rect 102002 10446 102004 10498
rect 101948 10386 102004 10446
rect 101948 10334 101950 10386
rect 102002 10334 102004 10386
rect 101948 10322 102004 10334
rect 102284 10498 102452 10500
rect 102284 10446 102398 10498
rect 102450 10446 102452 10498
rect 102284 10444 102452 10446
rect 101836 8318 101838 8370
rect 101890 8318 101892 8370
rect 101836 8306 101892 8318
rect 101948 8146 102004 8158
rect 101948 8094 101950 8146
rect 102002 8094 102004 8146
rect 101276 5854 101278 5906
rect 101330 5854 101332 5906
rect 101276 5842 101332 5854
rect 101388 6524 101780 6580
rect 101836 7586 101892 7598
rect 101836 7534 101838 7586
rect 101890 7534 101892 7586
rect 101836 6580 101892 7534
rect 101948 6692 102004 8094
rect 101948 6636 102228 6692
rect 101052 4562 101220 4564
rect 101052 4510 101054 4562
rect 101106 4510 101220 4562
rect 101052 4508 101220 4510
rect 101276 4900 101332 4910
rect 101052 4498 101108 4508
rect 101164 4340 101220 4350
rect 101276 4340 101332 4844
rect 101164 4338 101332 4340
rect 101164 4286 101166 4338
rect 101218 4286 101332 4338
rect 101164 4284 101332 4286
rect 101164 4274 101220 4284
rect 101388 4228 101444 6524
rect 101836 6514 101892 6524
rect 101612 6356 101668 6366
rect 102172 6356 102228 6636
rect 101500 5682 101556 5694
rect 101500 5630 101502 5682
rect 101554 5630 101556 5682
rect 101500 4452 101556 5630
rect 101612 5122 101668 6300
rect 101948 6300 102228 6356
rect 102284 6356 102340 10444
rect 102396 10434 102452 10444
rect 102508 11284 102564 11294
rect 102396 9716 102452 9726
rect 102508 9716 102564 11228
rect 102844 11172 102900 11182
rect 103404 11172 103460 11342
rect 104188 11284 104244 11294
rect 104188 11282 104356 11284
rect 104188 11230 104190 11282
rect 104242 11230 104356 11282
rect 104188 11228 104356 11230
rect 104188 11218 104244 11228
rect 102844 11170 103460 11172
rect 102844 11118 102846 11170
rect 102898 11118 103460 11170
rect 102844 11116 103460 11118
rect 102732 10276 102788 10286
rect 102732 9826 102788 10220
rect 102732 9774 102734 9826
rect 102786 9774 102788 9826
rect 102732 9762 102788 9774
rect 102396 9714 102564 9716
rect 102396 9662 102398 9714
rect 102450 9662 102564 9714
rect 102396 9660 102564 9662
rect 102396 9650 102452 9660
rect 102844 9044 102900 11116
rect 103628 10836 103684 10846
rect 103516 10724 103572 10734
rect 103516 10630 103572 10668
rect 102844 8978 102900 8988
rect 102956 10500 103012 10510
rect 102396 8484 102452 8494
rect 102956 8484 103012 10444
rect 103292 10276 103348 10286
rect 102396 8260 102452 8428
rect 102732 8428 103012 8484
rect 103068 10164 103124 10174
rect 102396 8204 102564 8260
rect 102396 8036 102452 8046
rect 102396 7942 102452 7980
rect 102508 7812 102564 8204
rect 102396 7756 102564 7812
rect 102732 7812 102788 8428
rect 103068 8372 103124 10108
rect 103292 9938 103348 10220
rect 103292 9886 103294 9938
rect 103346 9886 103348 9938
rect 103292 9874 103348 9886
rect 103628 9940 103684 10780
rect 104300 10834 104356 11228
rect 104300 10782 104302 10834
rect 104354 10782 104356 10834
rect 104300 10770 104356 10782
rect 104188 10724 104244 10734
rect 104188 10630 104244 10668
rect 104412 10612 104468 25452
rect 106092 23828 106148 116172
rect 106316 115890 106372 116396
rect 107660 116452 107716 116462
rect 107660 116358 107716 116396
rect 106316 115838 106318 115890
rect 106370 115838 106372 115890
rect 106316 115826 106372 115838
rect 107996 115780 108052 119200
rect 111132 117010 111188 119200
rect 111132 116958 111134 117010
rect 111186 116958 111188 117010
rect 111132 116946 111188 116958
rect 112252 117010 112308 117022
rect 112252 116958 112254 117010
rect 112306 116958 112308 117010
rect 108332 116564 108388 116574
rect 108332 116470 108388 116508
rect 112252 116562 112308 116958
rect 112700 117010 112756 119200
rect 112700 116958 112702 117010
rect 112754 116958 112756 117010
rect 112700 116946 112756 116958
rect 113596 117010 113652 117022
rect 113596 116958 113598 117010
rect 113650 116958 113652 117010
rect 112252 116510 112254 116562
rect 112306 116510 112308 116562
rect 112252 116498 112308 116510
rect 113596 116562 113652 116958
rect 115836 116676 115892 119200
rect 115836 116610 115892 116620
rect 116732 116676 116788 116686
rect 113596 116510 113598 116562
rect 113650 116510 113652 116562
rect 113596 116498 113652 116510
rect 116732 116562 116788 116620
rect 116732 116510 116734 116562
rect 116786 116510 116788 116562
rect 116732 116498 116788 116510
rect 111580 116452 111636 116462
rect 111132 116450 111636 116452
rect 111132 116398 111582 116450
rect 111634 116398 111636 116450
rect 111132 116396 111636 116398
rect 111132 115890 111188 116396
rect 111580 116386 111636 116396
rect 114380 116450 114436 116462
rect 116060 116452 116116 116462
rect 114380 116398 114382 116450
rect 114434 116398 114436 116450
rect 111996 116060 112260 116070
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 111996 115994 112260 116004
rect 111132 115838 111134 115890
rect 111186 115838 111188 115890
rect 111132 115826 111188 115838
rect 107996 115714 108052 115724
rect 108556 115780 108612 115790
rect 108556 115686 108612 115724
rect 109228 115666 109284 115678
rect 109228 115614 109230 115666
rect 109282 115614 109284 115666
rect 109228 115556 109284 115614
rect 110460 115668 110516 115678
rect 110012 115556 110068 115566
rect 109228 115554 110068 115556
rect 109228 115502 110014 115554
rect 110066 115502 110068 115554
rect 109228 115500 110068 115502
rect 105756 14644 105812 14654
rect 105196 12178 105252 12190
rect 105196 12126 105198 12178
rect 105250 12126 105252 12178
rect 104300 10556 104468 10612
rect 104524 12068 104580 12078
rect 105196 12068 105252 12126
rect 104524 12066 105252 12068
rect 104524 12014 104526 12066
rect 104578 12014 105252 12066
rect 104524 12012 105252 12014
rect 105420 12068 105476 12078
rect 104076 10388 104132 10398
rect 103964 10276 104020 10286
rect 103628 9938 103796 9940
rect 103628 9886 103630 9938
rect 103682 9886 103796 9938
rect 103628 9884 103796 9886
rect 103628 9874 103684 9884
rect 103628 8932 103684 8942
rect 102844 8316 103124 8372
rect 103404 8930 103684 8932
rect 103404 8878 103630 8930
rect 103682 8878 103684 8930
rect 103404 8876 103684 8878
rect 102844 8258 102900 8316
rect 102844 8206 102846 8258
rect 102898 8206 102900 8258
rect 102844 8194 102900 8206
rect 102956 7924 103012 7934
rect 102732 7756 102900 7812
rect 102396 7698 102452 7756
rect 102396 7646 102398 7698
rect 102450 7646 102452 7698
rect 102396 7252 102452 7646
rect 102732 7476 102788 7486
rect 102732 7382 102788 7420
rect 102396 7196 102788 7252
rect 101724 6130 101780 6142
rect 101724 6078 101726 6130
rect 101778 6078 101780 6130
rect 101724 5348 101780 6078
rect 101836 6020 101892 6030
rect 101836 5926 101892 5964
rect 101724 5282 101780 5292
rect 101612 5070 101614 5122
rect 101666 5070 101668 5122
rect 101612 5058 101668 5070
rect 101500 4386 101556 4396
rect 101836 5010 101892 5022
rect 101836 4958 101838 5010
rect 101890 4958 101892 5010
rect 101724 4340 101780 4350
rect 101612 4338 101780 4340
rect 101612 4286 101726 4338
rect 101778 4286 101780 4338
rect 101612 4284 101780 4286
rect 101612 4228 101668 4284
rect 101724 4274 101780 4284
rect 101836 4340 101892 4958
rect 101948 4564 102004 6300
rect 102284 6290 102340 6300
rect 102396 7028 102452 7038
rect 102060 5906 102116 5918
rect 102060 5854 102062 5906
rect 102114 5854 102116 5906
rect 102060 5572 102116 5854
rect 102396 5572 102452 6972
rect 102060 5516 102228 5572
rect 102060 5348 102116 5358
rect 102060 5254 102116 5292
rect 102060 4564 102116 4574
rect 101948 4562 102116 4564
rect 101948 4510 102062 4562
rect 102114 4510 102116 4562
rect 101948 4508 102116 4510
rect 102060 4498 102116 4508
rect 102172 4564 102228 5516
rect 102284 5516 102452 5572
rect 102508 6804 102564 6814
rect 102284 5234 102340 5516
rect 102284 5182 102286 5234
rect 102338 5182 102340 5234
rect 102284 5170 102340 5182
rect 102396 5348 102452 5358
rect 102396 5010 102452 5292
rect 102508 5122 102564 6748
rect 102732 6802 102788 7196
rect 102732 6750 102734 6802
rect 102786 6750 102788 6802
rect 102732 6738 102788 6750
rect 102620 6690 102676 6702
rect 102620 6638 102622 6690
rect 102674 6638 102676 6690
rect 102620 6580 102676 6638
rect 102620 6514 102676 6524
rect 102508 5070 102510 5122
rect 102562 5070 102564 5122
rect 102508 5058 102564 5070
rect 102396 4958 102398 5010
rect 102450 4958 102452 5010
rect 102396 4946 102452 4958
rect 102844 5012 102900 7756
rect 102844 4946 102900 4956
rect 102956 6018 103012 7868
rect 103404 7698 103460 8876
rect 103628 8866 103684 8876
rect 103740 8258 103796 9884
rect 103740 8206 103742 8258
rect 103794 8206 103796 8258
rect 103740 8194 103796 8206
rect 103964 8146 104020 10220
rect 103964 8094 103966 8146
rect 104018 8094 104020 8146
rect 103964 8082 104020 8094
rect 104076 9938 104132 10332
rect 104076 9886 104078 9938
rect 104130 9886 104132 9938
rect 103404 7646 103406 7698
rect 103458 7646 103460 7698
rect 103404 7634 103460 7646
rect 103516 8036 103572 8046
rect 103516 7698 103572 7980
rect 103516 7646 103518 7698
rect 103570 7646 103572 7698
rect 103516 7634 103572 7646
rect 103628 7476 103684 7486
rect 103292 7250 103348 7262
rect 103292 7198 103294 7250
rect 103346 7198 103348 7250
rect 103068 6580 103124 6590
rect 103068 6578 103236 6580
rect 103068 6526 103070 6578
rect 103122 6526 103236 6578
rect 103068 6524 103236 6526
rect 103068 6514 103124 6524
rect 103068 6356 103124 6366
rect 103068 6130 103124 6300
rect 103068 6078 103070 6130
rect 103122 6078 103124 6130
rect 103068 6066 103124 6078
rect 102956 5966 102958 6018
rect 103010 5966 103012 6018
rect 102956 4900 103012 5966
rect 103068 5682 103124 5694
rect 103068 5630 103070 5682
rect 103122 5630 103124 5682
rect 103068 5010 103124 5630
rect 103180 5124 103236 6524
rect 103292 5348 103348 7198
rect 103292 5282 103348 5292
rect 103180 5068 103348 5124
rect 103068 4958 103070 5010
rect 103122 4958 103124 5010
rect 103068 4946 103124 4958
rect 102956 4834 103012 4844
rect 103292 4900 103348 5068
rect 103292 4834 103348 4844
rect 103628 4898 103684 7420
rect 104076 7140 104132 9886
rect 104300 9268 104356 10556
rect 104412 10386 104468 10398
rect 104412 10334 104414 10386
rect 104466 10334 104468 10386
rect 104412 10050 104468 10334
rect 104412 9998 104414 10050
rect 104466 9998 104468 10050
rect 104412 9986 104468 9998
rect 104188 9212 104356 9268
rect 104188 8372 104244 9212
rect 104300 9044 104356 9054
rect 104300 8950 104356 8988
rect 104524 8932 104580 12012
rect 104748 11508 104804 11518
rect 104524 8866 104580 8876
rect 104636 10050 104692 10062
rect 104636 9998 104638 10050
rect 104690 9998 104692 10050
rect 104636 9602 104692 9998
rect 104636 9550 104638 9602
rect 104690 9550 104692 9602
rect 104188 8316 104356 8372
rect 104300 7698 104356 8316
rect 104412 8260 104468 8270
rect 104412 8166 104468 8204
rect 104300 7646 104302 7698
rect 104354 7646 104356 7698
rect 104188 7588 104244 7598
rect 104188 7494 104244 7532
rect 104300 7364 104356 7646
rect 103852 7084 104132 7140
rect 104188 7308 104356 7364
rect 104188 7252 104244 7308
rect 103852 6356 103908 7084
rect 103964 6916 104020 6926
rect 104188 6916 104244 7196
rect 104636 7028 104692 9550
rect 103964 6690 104020 6860
rect 103964 6638 103966 6690
rect 104018 6638 104020 6690
rect 103964 6626 104020 6638
rect 104076 6860 104244 6916
rect 104300 6972 104692 7028
rect 104076 6468 104132 6860
rect 104188 6692 104244 6702
rect 104188 6598 104244 6636
rect 104076 6412 104244 6468
rect 103908 6300 104132 6356
rect 103852 6290 103908 6300
rect 104076 6018 104132 6300
rect 104076 5966 104078 6018
rect 104130 5966 104132 6018
rect 104076 5572 104132 5966
rect 104076 5506 104132 5516
rect 103740 5124 103796 5134
rect 103740 5030 103796 5068
rect 104188 5122 104244 6412
rect 104188 5070 104190 5122
rect 104242 5070 104244 5122
rect 104188 5058 104244 5070
rect 103628 4846 103630 4898
rect 103682 4846 103684 4898
rect 103628 4834 103684 4846
rect 102172 4498 102228 4508
rect 102956 4450 103012 4462
rect 102956 4398 102958 4450
rect 103010 4398 103012 4450
rect 101948 4340 102004 4350
rect 101836 4338 102004 4340
rect 101836 4286 101950 4338
rect 102002 4286 102004 4338
rect 101836 4284 102004 4286
rect 101388 4172 101668 4228
rect 100716 3444 100772 3482
rect 100716 3378 100772 3388
rect 101164 3444 101220 3454
rect 100492 1362 100548 1372
rect 101164 800 101220 3388
rect 101836 3332 101892 4284
rect 101948 4274 102004 4284
rect 102172 4340 102228 4350
rect 102172 4246 102228 4284
rect 102396 4338 102452 4350
rect 102396 4286 102398 4338
rect 102450 4286 102452 4338
rect 102396 3780 102452 4286
rect 102396 3714 102452 3724
rect 102844 3556 102900 3566
rect 102956 3556 103012 4398
rect 103292 4452 103348 4462
rect 103292 4358 103348 4396
rect 104188 4340 104244 4350
rect 104188 4246 104244 4284
rect 104300 3892 104356 6972
rect 104412 6692 104468 6702
rect 104412 6356 104468 6636
rect 104524 6580 104580 6590
rect 104524 6486 104580 6524
rect 104412 6244 104468 6300
rect 104412 6188 104580 6244
rect 104412 6018 104468 6030
rect 104412 5966 104414 6018
rect 104466 5966 104468 6018
rect 104412 5012 104468 5966
rect 104412 4946 104468 4956
rect 104524 4788 104580 6188
rect 104524 4722 104580 4732
rect 104748 5010 104804 11452
rect 105420 10834 105476 12012
rect 105756 10836 105812 14588
rect 105980 12068 106036 12078
rect 105980 11974 106036 12012
rect 105420 10782 105422 10834
rect 105474 10782 105476 10834
rect 105420 10770 105476 10782
rect 105644 10780 105756 10836
rect 105308 10724 105364 10734
rect 105196 9940 105252 9950
rect 105308 9940 105364 10668
rect 105532 10386 105588 10398
rect 105532 10334 105534 10386
rect 105586 10334 105588 10386
rect 105532 10164 105588 10334
rect 105532 10098 105588 10108
rect 105644 9940 105700 10780
rect 105756 10770 105812 10780
rect 106092 10724 106148 23772
rect 108668 27188 108724 27198
rect 108668 20188 108724 27132
rect 108668 20132 108836 20188
rect 107100 18564 107156 18574
rect 106876 14084 106932 14094
rect 106764 12068 106820 12078
rect 106652 11394 106708 11406
rect 106652 11342 106654 11394
rect 106706 11342 106708 11394
rect 106428 11172 106484 11182
rect 106428 11170 106596 11172
rect 106428 11118 106430 11170
rect 106482 11118 106596 11170
rect 106428 11116 106596 11118
rect 106428 11106 106484 11116
rect 106428 10836 106484 10846
rect 106428 10742 106484 10780
rect 105196 9938 105364 9940
rect 105196 9886 105198 9938
rect 105250 9886 105364 9938
rect 105196 9884 105364 9886
rect 105420 9884 105700 9940
rect 105980 10668 106148 10724
rect 105196 9874 105252 9884
rect 105196 9042 105252 9054
rect 105196 8990 105198 9042
rect 105250 8990 105252 9042
rect 105196 8932 105252 8990
rect 105196 8866 105252 8876
rect 105196 8596 105252 8606
rect 105196 8370 105252 8540
rect 105196 8318 105198 8370
rect 105250 8318 105252 8370
rect 105196 8306 105252 8318
rect 104860 8260 104916 8270
rect 104860 5684 104916 8204
rect 105308 8146 105364 8158
rect 105308 8094 105310 8146
rect 105362 8094 105364 8146
rect 105084 8036 105140 8046
rect 105084 7942 105140 7980
rect 105084 7364 105140 7374
rect 104972 7362 105140 7364
rect 104972 7310 105086 7362
rect 105138 7310 105140 7362
rect 104972 7308 105140 7310
rect 104972 5908 105028 7308
rect 105084 7298 105140 7308
rect 105084 6692 105140 6702
rect 105084 6598 105140 6636
rect 105308 6692 105364 8094
rect 105308 6626 105364 6636
rect 105420 6356 105476 9884
rect 105532 9602 105588 9614
rect 105532 9550 105534 9602
rect 105586 9550 105588 9602
rect 105532 8932 105588 9550
rect 105980 9604 106036 10668
rect 106092 10498 106148 10510
rect 106092 10446 106094 10498
rect 106146 10446 106148 10498
rect 106092 10164 106148 10446
rect 106092 10098 106148 10108
rect 106428 10388 106484 10398
rect 106428 9938 106484 10332
rect 106540 10386 106596 11116
rect 106540 10334 106542 10386
rect 106594 10334 106596 10386
rect 106540 10322 106596 10334
rect 106652 10388 106708 11342
rect 106652 10322 106708 10332
rect 106428 9886 106430 9938
rect 106482 9886 106484 9938
rect 106428 9874 106484 9886
rect 106540 10050 106596 10062
rect 106540 9998 106542 10050
rect 106594 9998 106596 10050
rect 106036 9548 106148 9604
rect 105980 9510 106036 9548
rect 105532 8260 105588 8876
rect 105980 8930 106036 8942
rect 105980 8878 105982 8930
rect 106034 8878 106036 8930
rect 105532 8194 105588 8204
rect 105644 8820 105700 8830
rect 105532 7700 105588 7710
rect 105644 7700 105700 8764
rect 105980 8596 106036 8878
rect 105980 8530 106036 8540
rect 106092 8484 106148 9548
rect 106092 8418 106148 8428
rect 105756 8036 105812 8046
rect 105756 7942 105812 7980
rect 106204 8034 106260 8046
rect 106204 7982 106206 8034
rect 106258 7982 106260 8034
rect 105588 7644 105700 7700
rect 105532 7568 105588 7644
rect 105756 7588 105812 7598
rect 105644 6580 105700 6590
rect 105644 6486 105700 6524
rect 104972 5842 105028 5852
rect 105308 6300 105476 6356
rect 104860 5628 105140 5684
rect 104748 4958 104750 5010
rect 104802 4958 104804 5010
rect 104412 4450 104468 4462
rect 104412 4398 104414 4450
rect 104466 4398 104468 4450
rect 104412 4004 104468 4398
rect 104748 4452 104804 4958
rect 104748 4386 104804 4396
rect 104412 3948 104916 4004
rect 104300 3836 104692 3892
rect 102844 3554 103012 3556
rect 102844 3502 102846 3554
rect 102898 3502 103012 3554
rect 102844 3500 103012 3502
rect 102844 3490 102900 3500
rect 101948 3444 102004 3482
rect 101948 3378 102004 3388
rect 104076 3444 104132 3482
rect 104076 3378 104132 3388
rect 104524 3444 104580 3454
rect 101836 3266 101892 3276
rect 102844 3332 102900 3342
rect 102844 800 102900 3276
rect 104524 800 104580 3388
rect 104636 3332 104692 3836
rect 104748 3668 104804 3678
rect 104860 3668 104916 3948
rect 104972 3668 105028 3678
rect 104860 3666 105028 3668
rect 104860 3614 104974 3666
rect 105026 3614 105028 3666
rect 104860 3612 105028 3614
rect 104748 3554 104804 3612
rect 104972 3602 105028 3612
rect 104748 3502 104750 3554
rect 104802 3502 104804 3554
rect 104748 3490 104804 3502
rect 104636 3266 104692 3276
rect 105084 2212 105140 5628
rect 105196 5572 105252 5582
rect 105196 4116 105252 5516
rect 105308 5122 105364 6300
rect 105644 6132 105700 6142
rect 105644 5906 105700 6076
rect 105644 5854 105646 5906
rect 105698 5854 105700 5906
rect 105644 5842 105700 5854
rect 105420 5796 105476 5806
rect 105420 5702 105476 5740
rect 105644 5684 105700 5694
rect 105644 5348 105700 5628
rect 105308 5070 105310 5122
rect 105362 5070 105364 5122
rect 105308 5058 105364 5070
rect 105420 5236 105476 5246
rect 105308 4788 105364 4798
rect 105420 4788 105476 5180
rect 105644 5122 105700 5292
rect 105644 5070 105646 5122
rect 105698 5070 105700 5122
rect 105644 5058 105700 5070
rect 105532 4898 105588 4910
rect 105532 4846 105534 4898
rect 105586 4846 105588 4898
rect 105532 4788 105588 4846
rect 105364 4732 105588 4788
rect 105308 4722 105364 4732
rect 105756 4676 105812 7532
rect 106204 7588 106260 7982
rect 106204 7522 106260 7532
rect 106428 7476 106484 7486
rect 106428 7382 106484 7420
rect 105980 7362 106036 7374
rect 105980 7310 105982 7362
rect 106034 7310 106036 7362
rect 105868 6802 105924 6814
rect 105868 6750 105870 6802
rect 105922 6750 105924 6802
rect 105868 6580 105924 6750
rect 105868 5124 105924 6524
rect 105980 6468 106036 7310
rect 105980 6402 106036 6412
rect 106092 6692 106148 6702
rect 105868 5058 105924 5068
rect 105980 5010 106036 5022
rect 105980 4958 105982 5010
rect 106034 4958 106036 5010
rect 105980 4900 106036 4958
rect 105980 4834 106036 4844
rect 106092 4898 106148 6636
rect 106316 5796 106372 5806
rect 106540 5796 106596 9998
rect 106652 8036 106708 8046
rect 106652 7942 106708 7980
rect 106316 5794 106484 5796
rect 106316 5742 106318 5794
rect 106370 5742 106484 5794
rect 106316 5740 106484 5742
rect 106316 5730 106372 5740
rect 106316 5236 106372 5246
rect 106316 5142 106372 5180
rect 106092 4846 106094 4898
rect 106146 4846 106148 4898
rect 106092 4834 106148 4846
rect 105420 4620 105812 4676
rect 105308 4564 105364 4574
rect 105308 4470 105364 4508
rect 105420 4562 105476 4620
rect 105420 4510 105422 4562
rect 105474 4510 105476 4562
rect 105420 4340 105476 4510
rect 106428 4564 106484 5740
rect 106540 5730 106596 5740
rect 106652 7140 106708 7150
rect 106652 6578 106708 7084
rect 106764 6916 106820 12012
rect 106876 8148 106932 14028
rect 107100 11170 107156 18508
rect 107100 11118 107102 11170
rect 107154 11118 107156 11170
rect 106988 10498 107044 10510
rect 106988 10446 106990 10498
rect 107042 10446 107044 10498
rect 106988 10388 107044 10446
rect 106988 10322 107044 10332
rect 106988 10050 107044 10062
rect 106988 9998 106990 10050
rect 107042 9998 107044 10050
rect 106988 9938 107044 9998
rect 106988 9886 106990 9938
rect 107042 9886 107044 9938
rect 106988 9874 107044 9886
rect 107100 9716 107156 11118
rect 106876 8082 106932 8092
rect 106988 9660 107156 9716
rect 107212 12740 107268 12750
rect 106876 7924 106932 7934
rect 106876 7698 106932 7868
rect 106876 7646 106878 7698
rect 106930 7646 106932 7698
rect 106876 7634 106932 7646
rect 106764 6860 106932 6916
rect 106764 6692 106820 6702
rect 106764 6598 106820 6636
rect 106652 6526 106654 6578
rect 106706 6526 106708 6578
rect 106652 5460 106708 6526
rect 106652 5394 106708 5404
rect 106876 6132 106932 6860
rect 106876 6018 106932 6076
rect 106876 5966 106878 6018
rect 106930 5966 106932 6018
rect 106764 5346 106820 5358
rect 106764 5294 106766 5346
rect 106818 5294 106820 5346
rect 106652 5236 106708 5246
rect 106764 5236 106820 5294
rect 106652 5234 106820 5236
rect 106652 5182 106654 5234
rect 106706 5182 106820 5234
rect 106652 5180 106820 5182
rect 106652 5170 106708 5180
rect 106428 4498 106484 4508
rect 106540 5012 106596 5022
rect 105420 4274 105476 4284
rect 105644 4338 105700 4350
rect 105644 4286 105646 4338
rect 105698 4286 105700 4338
rect 105644 4116 105700 4286
rect 105980 4340 106036 4350
rect 105980 4246 106036 4284
rect 106540 4338 106596 4956
rect 106540 4286 106542 4338
rect 106594 4286 106596 4338
rect 106540 4274 106596 4286
rect 105196 4060 105700 4116
rect 106204 4228 106260 4238
rect 105532 3666 105588 3678
rect 105532 3614 105534 3666
rect 105586 3614 105588 3666
rect 105532 3554 105588 3614
rect 105532 3502 105534 3554
rect 105586 3502 105588 3554
rect 105532 3490 105588 3502
rect 105084 2146 105140 2156
rect 106204 800 106260 4172
rect 106428 3444 106484 3482
rect 106428 3378 106484 3388
rect 106876 3220 106932 5966
rect 106988 5346 107044 9660
rect 107212 8484 107268 12684
rect 108668 12180 108724 12190
rect 108556 12178 108724 12180
rect 108556 12126 108670 12178
rect 108722 12126 108724 12178
rect 108556 12124 108724 12126
rect 108108 12068 108164 12078
rect 108108 11974 108164 12012
rect 107436 11618 107492 11630
rect 107436 11566 107438 11618
rect 107490 11566 107492 11618
rect 107436 11506 107492 11566
rect 107436 11454 107438 11506
rect 107490 11454 107492 11506
rect 107436 11442 107492 11454
rect 107884 11170 107940 11182
rect 108332 11172 108388 11182
rect 107884 11118 107886 11170
rect 107938 11118 107940 11170
rect 107884 10612 107940 11118
rect 107884 10546 107940 10556
rect 108108 11170 108388 11172
rect 108108 11118 108334 11170
rect 108386 11118 108388 11170
rect 108108 11116 108388 11118
rect 107100 8428 107268 8484
rect 107324 10498 107380 10510
rect 107324 10446 107326 10498
rect 107378 10446 107380 10498
rect 107324 10386 107380 10446
rect 107324 10334 107326 10386
rect 107378 10334 107380 10386
rect 107100 7700 107156 8428
rect 107100 7028 107156 7644
rect 107100 6962 107156 6972
rect 107212 8148 107268 8158
rect 107212 6804 107268 8092
rect 107212 6738 107268 6748
rect 107100 6692 107156 6702
rect 107100 6020 107156 6636
rect 107324 6692 107380 10334
rect 107436 9602 107492 9614
rect 107436 9550 107438 9602
rect 107490 9550 107492 9602
rect 107436 8484 107492 9550
rect 107884 9604 107940 9614
rect 108108 9604 108164 11116
rect 108332 10836 108388 11116
rect 108556 10836 108612 12124
rect 108668 12114 108724 12124
rect 108332 10834 108612 10836
rect 108332 10782 108558 10834
rect 108610 10782 108612 10834
rect 108332 10780 108612 10782
rect 108556 10770 108612 10780
rect 108332 10612 108388 10622
rect 107884 9602 108164 9604
rect 107884 9550 107886 9602
rect 107938 9550 108164 9602
rect 107884 9548 108164 9550
rect 108220 10498 108276 10510
rect 108220 10446 108222 10498
rect 108274 10446 108276 10498
rect 107884 9044 107940 9548
rect 107884 8978 107940 8988
rect 108108 8930 108164 8942
rect 108108 8878 108110 8930
rect 108162 8878 108164 8930
rect 108108 8820 108164 8878
rect 108108 8754 108164 8764
rect 107436 8428 107604 8484
rect 107436 7700 107492 7710
rect 107436 7606 107492 7644
rect 107324 6626 107380 6636
rect 107100 5926 107156 5964
rect 107436 6020 107492 6030
rect 107436 5906 107492 5964
rect 107436 5854 107438 5906
rect 107490 5854 107492 5906
rect 106988 5294 106990 5346
rect 107042 5294 107044 5346
rect 106988 5282 107044 5294
rect 107324 5794 107380 5806
rect 107324 5742 107326 5794
rect 107378 5742 107380 5794
rect 107324 4788 107380 5742
rect 107436 5796 107492 5854
rect 107436 5730 107492 5740
rect 107324 4722 107380 4732
rect 107548 4900 107604 8428
rect 107996 8036 108052 8046
rect 107996 7942 108052 7980
rect 107884 7924 107940 7934
rect 107660 7812 107716 7822
rect 107660 5572 107716 7756
rect 107660 5122 107716 5516
rect 107772 7474 107828 7486
rect 107772 7422 107774 7474
rect 107826 7422 107828 7474
rect 107772 5234 107828 7422
rect 107884 6020 107940 7868
rect 107996 7588 108052 7598
rect 107996 7028 108052 7532
rect 107996 6962 108052 6972
rect 108108 7588 108164 7598
rect 108220 7588 108276 10446
rect 108332 9938 108388 10556
rect 108668 10388 108724 10398
rect 108332 9886 108334 9938
rect 108386 9886 108388 9938
rect 108332 9874 108388 9886
rect 108556 10276 108612 10286
rect 108556 9268 108612 10220
rect 108332 9266 108612 9268
rect 108332 9214 108558 9266
rect 108610 9214 108612 9266
rect 108332 9212 108612 9214
rect 108332 8258 108388 9212
rect 108556 9202 108612 9212
rect 108668 9156 108724 10332
rect 108332 8206 108334 8258
rect 108386 8206 108388 8258
rect 108332 8194 108388 8206
rect 108444 8372 108500 8382
rect 108108 7586 108276 7588
rect 108108 7534 108110 7586
rect 108162 7534 108276 7586
rect 108108 7532 108276 7534
rect 107996 6020 108052 6030
rect 107884 6018 108052 6020
rect 107884 5966 107998 6018
rect 108050 5966 108052 6018
rect 107884 5964 108052 5966
rect 107996 5908 108052 5964
rect 107996 5842 108052 5852
rect 107772 5182 107774 5234
rect 107826 5182 107828 5234
rect 107772 5170 107828 5182
rect 107660 5070 107662 5122
rect 107714 5070 107716 5122
rect 107660 5058 107716 5070
rect 107100 4228 107156 4238
rect 107100 4134 107156 4172
rect 107548 4228 107604 4844
rect 108108 4340 108164 7532
rect 108220 7140 108276 7150
rect 108220 6356 108276 7084
rect 108220 6290 108276 6300
rect 108332 6020 108388 6030
rect 108108 4274 108164 4284
rect 108220 6018 108388 6020
rect 108220 5966 108334 6018
rect 108386 5966 108388 6018
rect 108220 5964 108388 5966
rect 107548 4162 107604 4172
rect 107548 3556 107604 3566
rect 107548 3462 107604 3500
rect 108220 3554 108276 5964
rect 108332 5954 108388 5964
rect 108332 5012 108388 5022
rect 108332 4918 108388 4956
rect 108332 4564 108388 4574
rect 108444 4564 108500 8316
rect 108556 7700 108612 7710
rect 108556 7362 108612 7644
rect 108556 7310 108558 7362
rect 108610 7310 108612 7362
rect 108556 6916 108612 7310
rect 108556 6850 108612 6860
rect 108332 4562 108500 4564
rect 108332 4510 108334 4562
rect 108386 4510 108500 4562
rect 108332 4508 108500 4510
rect 108556 5348 108612 5358
rect 108668 5348 108724 9100
rect 108780 8372 108836 20132
rect 109228 13636 109284 115500
rect 110012 115490 110068 115500
rect 110460 114994 110516 115612
rect 110796 115668 110852 115678
rect 110796 115574 110852 115612
rect 113036 115556 113092 115566
rect 113036 115462 113092 115500
rect 113932 115556 113988 115566
rect 110460 114942 110462 114994
rect 110514 114942 110516 114994
rect 110460 114930 110516 114942
rect 111996 114492 112260 114502
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 111996 114426 112260 114436
rect 111996 112924 112260 112934
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 111996 112858 112260 112868
rect 111996 111356 112260 111366
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 111996 111290 112260 111300
rect 111996 109788 112260 109798
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 111996 109722 112260 109732
rect 111996 108220 112260 108230
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 111996 108154 112260 108164
rect 111996 106652 112260 106662
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 111996 106586 112260 106596
rect 111996 105084 112260 105094
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 111996 105018 112260 105028
rect 111996 103516 112260 103526
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 111996 103450 112260 103460
rect 111996 101948 112260 101958
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 111996 101882 112260 101892
rect 111996 100380 112260 100390
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 111996 100314 112260 100324
rect 111996 98812 112260 98822
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 111996 98746 112260 98756
rect 111996 97244 112260 97254
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 111996 97178 112260 97188
rect 111996 95676 112260 95686
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 111996 95610 112260 95620
rect 111996 94108 112260 94118
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 111996 94042 112260 94052
rect 111996 92540 112260 92550
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 111996 92474 112260 92484
rect 111996 90972 112260 90982
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 111996 90906 112260 90916
rect 111996 89404 112260 89414
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 111996 89338 112260 89348
rect 111996 87836 112260 87846
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 111996 87770 112260 87780
rect 111996 86268 112260 86278
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 111996 86202 112260 86212
rect 111996 84700 112260 84710
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 111996 84634 112260 84644
rect 111996 83132 112260 83142
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 111996 83066 112260 83076
rect 111996 81564 112260 81574
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 111996 81498 112260 81508
rect 111996 79996 112260 80006
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 111996 79930 112260 79940
rect 111996 78428 112260 78438
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 111996 78362 112260 78372
rect 111996 76860 112260 76870
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 111996 76794 112260 76804
rect 111996 75292 112260 75302
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 111996 75226 112260 75236
rect 111996 73724 112260 73734
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 111996 73658 112260 73668
rect 111996 72156 112260 72166
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 111996 72090 112260 72100
rect 111996 70588 112260 70598
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 111996 70522 112260 70532
rect 111996 69020 112260 69030
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 111996 68954 112260 68964
rect 111996 67452 112260 67462
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 111996 67386 112260 67396
rect 111996 65884 112260 65894
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 111996 65818 112260 65828
rect 111996 64316 112260 64326
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 111996 64250 112260 64260
rect 111996 62748 112260 62758
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 111996 62682 112260 62692
rect 111996 61180 112260 61190
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 111996 61114 112260 61124
rect 111996 59612 112260 59622
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 111996 59546 112260 59556
rect 111996 58044 112260 58054
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 111996 57978 112260 57988
rect 111996 56476 112260 56486
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 111996 56410 112260 56420
rect 111996 54908 112260 54918
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 111996 54842 112260 54852
rect 111996 53340 112260 53350
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 111996 53274 112260 53284
rect 111996 51772 112260 51782
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 111996 51706 112260 51716
rect 111996 50204 112260 50214
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 111996 50138 112260 50148
rect 111996 48636 112260 48646
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 111996 48570 112260 48580
rect 111996 47068 112260 47078
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 111996 47002 112260 47012
rect 111996 45500 112260 45510
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 111996 45434 112260 45444
rect 111996 43932 112260 43942
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 111996 43866 112260 43876
rect 111996 42364 112260 42374
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 111996 42298 112260 42308
rect 111996 40796 112260 40806
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 111996 40730 112260 40740
rect 111996 39228 112260 39238
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 111996 39162 112260 39172
rect 111996 37660 112260 37670
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 111996 37594 112260 37604
rect 111996 36092 112260 36102
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 111996 36026 112260 36036
rect 111996 34524 112260 34534
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 111996 34458 112260 34468
rect 111996 32956 112260 32966
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 111996 32890 112260 32900
rect 111996 31388 112260 31398
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 111996 31322 112260 31332
rect 111996 29820 112260 29830
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 111996 29754 112260 29764
rect 111996 28252 112260 28262
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 111996 28186 112260 28196
rect 111996 26684 112260 26694
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 111996 26618 112260 26628
rect 111996 25116 112260 25126
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 111996 25050 112260 25060
rect 112364 23716 112420 23726
rect 111996 23548 112260 23558
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 111996 23482 112260 23492
rect 111996 21980 112260 21990
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 111996 21914 112260 21924
rect 111996 20412 112260 20422
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 111996 20346 112260 20356
rect 111996 18844 112260 18854
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 111996 18778 112260 18788
rect 111996 17276 112260 17286
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 111996 17210 112260 17220
rect 111996 15708 112260 15718
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 111996 15642 112260 15652
rect 111996 14140 112260 14150
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 111996 14074 112260 14084
rect 109228 13570 109284 13580
rect 111580 13636 111636 13646
rect 109452 12068 109508 12078
rect 109452 11974 109508 12012
rect 111580 12066 111636 13580
rect 111996 12572 112260 12582
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 111996 12506 112260 12516
rect 111580 12014 111582 12066
rect 111634 12014 111636 12066
rect 110796 11844 110852 11854
rect 109116 11396 109172 11406
rect 109004 11394 109284 11396
rect 109004 11342 109118 11394
rect 109170 11342 109284 11394
rect 109004 11340 109284 11342
rect 109004 10612 109060 11340
rect 109116 11330 109172 11340
rect 109004 10546 109060 10556
rect 109116 10610 109172 10622
rect 109116 10558 109118 10610
rect 109170 10558 109172 10610
rect 109116 9044 109172 10558
rect 109228 9826 109284 11340
rect 109900 11282 109956 11294
rect 109900 11230 109902 11282
rect 109954 11230 109956 11282
rect 109900 11172 109956 11230
rect 109900 11106 109956 11116
rect 110460 10836 110516 10846
rect 109900 10498 109956 10510
rect 109900 10446 109902 10498
rect 109954 10446 109956 10498
rect 109900 10276 109956 10446
rect 109900 10210 109956 10220
rect 109228 9774 109230 9826
rect 109282 9774 109284 9826
rect 109228 9762 109284 9774
rect 110012 9714 110068 9726
rect 110012 9662 110014 9714
rect 110066 9662 110068 9714
rect 110012 9604 110068 9662
rect 110012 9538 110068 9548
rect 109116 8950 109172 8988
rect 110012 9044 110068 9054
rect 109900 8932 109956 8942
rect 109900 8838 109956 8876
rect 109676 8708 109732 8718
rect 108780 8306 108836 8316
rect 109564 8596 109620 8606
rect 109340 8260 109396 8270
rect 109396 8204 109508 8260
rect 109340 8128 109396 8204
rect 109228 8036 109284 8046
rect 109004 7362 109060 7374
rect 109004 7310 109006 7362
rect 109058 7310 109060 7362
rect 109004 7140 109060 7310
rect 109004 7074 109060 7084
rect 108612 5292 108724 5348
rect 109116 6578 109172 6590
rect 109116 6526 109118 6578
rect 109170 6526 109172 6578
rect 108332 4498 108388 4508
rect 108444 4338 108500 4350
rect 108444 4286 108446 4338
rect 108498 4286 108500 4338
rect 108444 4228 108500 4286
rect 108556 4338 108612 5292
rect 109116 5236 109172 6526
rect 109228 6468 109284 7980
rect 109340 7250 109396 7262
rect 109340 7198 109342 7250
rect 109394 7198 109396 7250
rect 109340 6802 109396 7198
rect 109340 6750 109342 6802
rect 109394 6750 109396 6802
rect 109340 6738 109396 6750
rect 109452 7252 109508 8204
rect 109564 7698 109620 8540
rect 109564 7646 109566 7698
rect 109618 7646 109620 7698
rect 109564 7634 109620 7646
rect 109340 6468 109396 6478
rect 109228 6412 109340 6468
rect 109340 6374 109396 6412
rect 109452 6244 109508 7196
rect 109228 6188 109508 6244
rect 109564 6468 109620 6478
rect 109228 5906 109284 6188
rect 109228 5854 109230 5906
rect 109282 5854 109284 5906
rect 109228 5842 109284 5854
rect 109452 5796 109508 5806
rect 109116 5180 109284 5236
rect 108892 5012 108948 5022
rect 108892 4450 108948 4956
rect 108892 4398 108894 4450
rect 108946 4398 108948 4450
rect 108892 4386 108948 4398
rect 109116 4898 109172 4910
rect 109116 4846 109118 4898
rect 109170 4846 109172 4898
rect 108556 4286 108558 4338
rect 108610 4286 108612 4338
rect 108556 4274 108612 4286
rect 108444 3892 108500 4172
rect 108444 3826 108500 3836
rect 109116 3668 109172 4846
rect 109228 4562 109284 5180
rect 109452 5122 109508 5740
rect 109452 5070 109454 5122
rect 109506 5070 109508 5122
rect 109452 5058 109508 5070
rect 109564 5124 109620 6412
rect 109564 5058 109620 5068
rect 109676 4788 109732 8652
rect 110012 8484 110068 8988
rect 110012 8372 110068 8428
rect 109900 8316 110068 8372
rect 110236 8820 110292 8830
rect 109900 7698 109956 8316
rect 109900 7646 109902 7698
rect 109954 7646 109956 7698
rect 109900 7634 109956 7646
rect 110012 8146 110068 8158
rect 110012 8094 110014 8146
rect 110066 8094 110068 8146
rect 110012 7250 110068 8094
rect 110012 7198 110014 7250
rect 110066 7198 110068 7250
rect 110012 7186 110068 7198
rect 110236 7700 110292 8764
rect 110236 6690 110292 7644
rect 110236 6638 110238 6690
rect 110290 6638 110292 6690
rect 110236 6626 110292 6638
rect 110348 7362 110404 7374
rect 110348 7310 110350 7362
rect 110402 7310 110404 7362
rect 110348 6580 110404 7310
rect 110348 6514 110404 6524
rect 110348 5908 110404 5918
rect 109900 5796 109956 5806
rect 109900 5794 110292 5796
rect 109900 5742 109902 5794
rect 109954 5742 110292 5794
rect 109900 5740 110292 5742
rect 109900 5730 109956 5740
rect 110236 5346 110292 5740
rect 110236 5294 110238 5346
rect 110290 5294 110292 5346
rect 110236 5282 110292 5294
rect 110236 5124 110292 5134
rect 110236 5030 110292 5068
rect 109228 4510 109230 4562
rect 109282 4510 109284 4562
rect 109228 4498 109284 4510
rect 109340 4732 109732 4788
rect 109228 4340 109284 4350
rect 109340 4340 109396 4732
rect 109228 4338 109396 4340
rect 109228 4286 109230 4338
rect 109282 4286 109396 4338
rect 109228 4284 109396 4286
rect 109900 4676 109956 4686
rect 109228 4274 109284 4284
rect 109452 4226 109508 4238
rect 109452 4174 109454 4226
rect 109506 4174 109508 4226
rect 109452 4116 109508 4174
rect 109452 4050 109508 4060
rect 109564 4228 109620 4238
rect 109116 3602 109172 3612
rect 108220 3502 108222 3554
rect 108274 3502 108276 3554
rect 108220 3490 108276 3502
rect 106876 3154 106932 3164
rect 107884 3444 107940 3454
rect 107884 800 107940 3388
rect 109004 3444 109060 3482
rect 109004 3378 109060 3388
rect 109564 800 109620 4172
rect 109900 3666 109956 4620
rect 110236 4228 110292 4238
rect 110236 4134 110292 4172
rect 109900 3614 109902 3666
rect 109954 3614 109956 3666
rect 109900 3602 109956 3614
rect 110348 3666 110404 5852
rect 110460 4676 110516 10780
rect 110796 8596 110852 11788
rect 111580 11844 111636 12014
rect 112140 12068 112196 12078
rect 112140 11974 112196 12012
rect 111580 11778 111636 11788
rect 112028 11508 112084 11518
rect 110796 8530 110852 8540
rect 111580 11506 112084 11508
rect 111580 11454 112030 11506
rect 112082 11454 112084 11506
rect 111580 11452 112084 11454
rect 111132 8036 111188 8046
rect 110796 7476 110852 7486
rect 110796 7382 110852 7420
rect 111132 6692 111188 7980
rect 111244 7362 111300 7374
rect 111244 7310 111246 7362
rect 111298 7310 111300 7362
rect 111244 7028 111300 7310
rect 111580 7364 111636 11452
rect 112028 11442 112084 11452
rect 111996 11004 112260 11014
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 111996 10938 112260 10948
rect 112028 10500 112084 10510
rect 112028 10164 112084 10444
rect 111692 10108 112084 10164
rect 111692 7812 111748 10108
rect 112140 10052 112196 10062
rect 111692 7746 111748 7756
rect 111804 9940 111860 9950
rect 111580 7298 111636 7308
rect 111244 6962 111300 6972
rect 111020 6690 111188 6692
rect 111020 6638 111134 6690
rect 111186 6638 111188 6690
rect 111020 6636 111188 6638
rect 110572 6468 110628 6478
rect 110572 6466 110740 6468
rect 110572 6414 110574 6466
rect 110626 6414 110740 6466
rect 110572 6412 110740 6414
rect 110572 6402 110628 6412
rect 110572 5010 110628 5022
rect 110572 4958 110574 5010
rect 110626 4958 110628 5010
rect 110572 4900 110628 4958
rect 110572 4834 110628 4844
rect 110460 4610 110516 4620
rect 110684 4340 110740 6412
rect 110796 6356 110852 6366
rect 110796 5908 110852 6300
rect 110796 5842 110852 5852
rect 111020 5796 111076 6636
rect 111132 6626 111188 6636
rect 111020 5730 111076 5740
rect 111132 6468 111188 6478
rect 111132 5572 111188 6412
rect 111244 6468 111300 6478
rect 111692 6468 111748 6478
rect 111244 6466 111748 6468
rect 111244 6414 111246 6466
rect 111298 6414 111694 6466
rect 111746 6414 111748 6466
rect 111244 6412 111748 6414
rect 111244 6402 111300 6412
rect 111132 5346 111188 5516
rect 111132 5294 111134 5346
rect 111186 5294 111188 5346
rect 111132 5282 111188 5294
rect 111356 5460 111412 6412
rect 111692 6402 111748 6412
rect 111356 4898 111412 5404
rect 111356 4846 111358 4898
rect 111410 4846 111412 4898
rect 111356 4452 111412 4846
rect 111356 4386 111412 4396
rect 111468 5348 111524 5358
rect 111020 4340 111076 4350
rect 110684 4338 111076 4340
rect 110684 4286 111022 4338
rect 111074 4286 111076 4338
rect 110684 4284 111076 4286
rect 111020 4274 111076 4284
rect 111468 4340 111524 5292
rect 111468 4274 111524 4284
rect 111804 4452 111860 9884
rect 112140 9938 112196 9996
rect 112140 9886 112142 9938
rect 112194 9886 112196 9938
rect 112140 9716 112196 9886
rect 112140 9650 112196 9660
rect 111996 9436 112260 9446
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 111996 9370 112260 9380
rect 112028 9044 112084 9054
rect 112028 8930 112084 8988
rect 112028 8878 112030 8930
rect 112082 8878 112084 8930
rect 112028 8866 112084 8878
rect 112252 8148 112308 8158
rect 112252 8034 112308 8092
rect 112252 7982 112254 8034
rect 112306 7982 112308 8034
rect 112252 7970 112308 7982
rect 111996 7868 112260 7878
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 111996 7802 112260 7812
rect 112364 7812 112420 23660
rect 113596 19348 113652 19358
rect 113260 16884 113316 16894
rect 112588 11844 112644 11854
rect 112588 8036 112644 11788
rect 112700 11170 112756 11182
rect 112700 11118 112702 11170
rect 112754 11118 112756 11170
rect 112700 11060 112756 11118
rect 113148 11172 113204 11182
rect 113148 11078 113204 11116
rect 112700 10994 112756 11004
rect 113148 10498 113204 10510
rect 113148 10446 113150 10498
rect 113202 10446 113204 10498
rect 113148 10276 113204 10446
rect 113148 10210 113204 10220
rect 113260 9940 113316 16828
rect 113596 15148 113652 19292
rect 113484 15092 113652 15148
rect 113484 10164 113540 15092
rect 113596 10500 113652 10510
rect 113596 10498 113764 10500
rect 113596 10446 113598 10498
rect 113650 10446 113764 10498
rect 113596 10444 113764 10446
rect 113596 10434 113652 10444
rect 113596 10164 113652 10174
rect 113484 10108 113596 10164
rect 113260 9938 113428 9940
rect 113260 9886 113262 9938
rect 113314 9886 113428 9938
rect 113260 9884 113428 9886
rect 113260 9874 113316 9884
rect 112812 9604 112868 9614
rect 112812 9510 112868 9548
rect 113036 9156 113092 9166
rect 113036 9062 113092 9100
rect 113260 8372 113316 8382
rect 113260 8278 113316 8316
rect 112588 7970 112644 7980
rect 112812 8034 112868 8046
rect 112812 7982 112814 8034
rect 112866 7982 112868 8034
rect 112364 7698 112420 7756
rect 112364 7646 112366 7698
rect 112418 7646 112420 7698
rect 112364 7634 112420 7646
rect 112812 7924 112868 7982
rect 112028 7474 112084 7486
rect 112028 7422 112030 7474
rect 112082 7422 112084 7474
rect 112028 7364 112084 7422
rect 112028 7298 112084 7308
rect 112812 7252 112868 7868
rect 113148 7588 113204 7598
rect 112812 7186 112868 7196
rect 112924 7586 113204 7588
rect 112924 7534 113150 7586
rect 113202 7534 113204 7586
rect 112924 7532 113204 7534
rect 112364 7028 112420 7038
rect 112140 6692 112196 6702
rect 112140 6598 112196 6636
rect 111996 6300 112260 6310
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 111996 6234 112260 6244
rect 112140 5796 112196 5806
rect 112364 5796 112420 6972
rect 112588 6466 112644 6478
rect 112588 6414 112590 6466
rect 112642 6414 112644 6466
rect 112588 6020 112644 6414
rect 112588 5954 112644 5964
rect 112140 5794 112420 5796
rect 112140 5742 112142 5794
rect 112194 5742 112420 5794
rect 112140 5740 112420 5742
rect 112140 5730 112196 5740
rect 112252 5348 112308 5358
rect 112252 5234 112308 5292
rect 112252 5182 112254 5234
rect 112306 5182 112308 5234
rect 112252 5170 112308 5182
rect 112364 5124 112420 5740
rect 112700 5908 112756 5918
rect 112588 5124 112644 5134
rect 112364 5122 112644 5124
rect 112364 5070 112590 5122
rect 112642 5070 112644 5122
rect 112364 5068 112644 5070
rect 112588 4788 112644 5068
rect 111996 4732 112260 4742
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112588 4722 112644 4732
rect 111996 4666 112260 4676
rect 112028 4452 112084 4462
rect 111804 4450 112084 4452
rect 111804 4398 112030 4450
rect 112082 4398 112084 4450
rect 111804 4396 112084 4398
rect 110348 3614 110350 3666
rect 110402 3614 110404 3666
rect 110348 3602 110404 3614
rect 110796 3780 110852 3790
rect 110796 3554 110852 3724
rect 110796 3502 110798 3554
rect 110850 3502 110852 3554
rect 110796 2324 110852 3502
rect 110796 2258 110852 2268
rect 111244 3444 111300 3454
rect 111244 800 111300 3388
rect 111804 1428 111860 4396
rect 112028 4386 112084 4396
rect 112364 4450 112420 4462
rect 112364 4398 112366 4450
rect 112418 4398 112420 4450
rect 112364 3556 112420 4398
rect 112364 3490 112420 3500
rect 111916 3444 111972 3482
rect 111916 3378 111972 3388
rect 111996 3164 112260 3174
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 111996 3098 112260 3108
rect 112700 2772 112756 5852
rect 112924 4564 112980 7532
rect 113148 7522 113204 7532
rect 113372 7474 113428 9884
rect 113372 7422 113374 7474
rect 113426 7422 113428 7474
rect 113372 7410 113428 7422
rect 113484 8930 113540 8942
rect 113484 8878 113486 8930
rect 113538 8878 113540 8930
rect 113484 7364 113540 8878
rect 113484 7298 113540 7308
rect 113036 6580 113092 6590
rect 113036 5236 113092 6524
rect 113484 6466 113540 6478
rect 113484 6414 113486 6466
rect 113538 6414 113540 6466
rect 113372 6244 113428 6254
rect 113148 5908 113204 5918
rect 113148 5814 113204 5852
rect 113372 5906 113428 6188
rect 113484 6132 113540 6414
rect 113484 6066 113540 6076
rect 113372 5854 113374 5906
rect 113426 5854 113428 5906
rect 113372 5842 113428 5854
rect 113596 5796 113652 10108
rect 113708 9602 113764 10444
rect 113932 10498 113988 115500
rect 114380 115556 114436 116398
rect 115836 116450 116116 116452
rect 115836 116398 116062 116450
rect 116114 116398 116116 116450
rect 115836 116396 116116 116398
rect 115836 115890 115892 116396
rect 116060 116386 116116 116396
rect 115836 115838 115838 115890
rect 115890 115838 115892 115890
rect 115836 115826 115892 115838
rect 117404 115780 117460 119200
rect 120540 116564 120596 119200
rect 120540 116498 120596 116508
rect 121436 116564 121492 116574
rect 121436 116470 121492 116508
rect 122108 116564 122164 119200
rect 125244 116676 125300 119200
rect 125244 116610 125300 116620
rect 126028 116676 126084 116686
rect 122108 116498 122164 116508
rect 124012 116564 124068 116574
rect 124012 116470 124068 116508
rect 126028 116562 126084 116620
rect 126028 116510 126030 116562
rect 126082 116510 126084 116562
rect 126028 116498 126084 116510
rect 126812 116564 126868 119200
rect 127356 116844 127620 116854
rect 127412 116788 127460 116844
rect 127516 116788 127564 116844
rect 127356 116778 127620 116788
rect 126812 116498 126868 116508
rect 127932 116564 127988 116574
rect 127932 116470 127988 116508
rect 129948 116564 130004 119200
rect 129948 116498 130004 116508
rect 120092 116452 120148 116462
rect 118972 116228 119028 116238
rect 117404 115714 117460 115724
rect 118524 115780 118580 115790
rect 118524 115686 118580 115724
rect 114940 115668 114996 115678
rect 114940 115574 114996 115612
rect 115500 115668 115556 115678
rect 115500 115574 115556 115612
rect 117628 115666 117684 115678
rect 117628 115614 117630 115666
rect 117682 115614 117684 115666
rect 114380 115490 114436 115500
rect 117180 115556 117236 115566
rect 117628 115556 117684 115614
rect 117180 115554 117684 115556
rect 117180 115502 117182 115554
rect 117234 115502 117684 115554
rect 117180 115500 117684 115502
rect 117180 102508 117236 115500
rect 116956 102452 117236 102508
rect 115052 20804 115108 20814
rect 114828 19796 114884 19806
rect 113932 10446 113934 10498
rect 113986 10446 113988 10498
rect 113932 9828 113988 10446
rect 114156 17668 114212 17678
rect 114156 9940 114212 17612
rect 114268 17108 114324 17118
rect 114268 10724 114324 17052
rect 114828 15148 114884 19740
rect 114828 15092 114996 15148
rect 114716 12404 114772 12414
rect 114716 11172 114772 12348
rect 114716 11078 114772 11116
rect 114268 10658 114324 10668
rect 114492 10500 114548 10510
rect 114380 10498 114548 10500
rect 114380 10446 114494 10498
rect 114546 10446 114548 10498
rect 114380 10444 114548 10446
rect 114268 10164 114324 10174
rect 114380 10164 114436 10444
rect 114492 10434 114548 10444
rect 114324 10108 114436 10164
rect 114268 10098 114324 10108
rect 114156 9808 114212 9884
rect 114828 10050 114884 10062
rect 114828 9998 114830 10050
rect 114882 9998 114884 10050
rect 113932 9762 113988 9772
rect 113708 9550 113710 9602
rect 113762 9550 113764 9602
rect 113708 9266 113764 9550
rect 114492 9716 114548 9726
rect 113708 9214 113710 9266
rect 113762 9214 113764 9266
rect 113708 9202 113764 9214
rect 114380 9268 114436 9278
rect 114380 9174 114436 9212
rect 114044 9044 114100 9054
rect 113708 9042 114100 9044
rect 113708 8990 114046 9042
rect 114098 8990 114100 9042
rect 113708 8988 114100 8990
rect 113708 8708 113764 8988
rect 114044 8978 114100 8988
rect 113708 8642 113764 8652
rect 113820 8818 113876 8830
rect 113820 8766 113822 8818
rect 113874 8766 113876 8818
rect 113708 8148 113764 8158
rect 113708 8054 113764 8092
rect 113820 7924 113876 8766
rect 113596 5702 113652 5740
rect 113708 7868 113876 7924
rect 114044 8708 114100 8718
rect 113708 5460 113764 7868
rect 113820 7364 113876 7374
rect 113820 6692 113876 7308
rect 113932 7362 113988 7374
rect 113932 7310 113934 7362
rect 113986 7310 113988 7362
rect 113932 7252 113988 7310
rect 113932 7186 113988 7196
rect 113932 6692 113988 6702
rect 113820 6690 113988 6692
rect 113820 6638 113934 6690
rect 113986 6638 113988 6690
rect 113820 6636 113988 6638
rect 113932 6626 113988 6636
rect 114044 6692 114100 8652
rect 114492 8484 114548 9660
rect 114716 9602 114772 9614
rect 114716 9550 114718 9602
rect 114770 9550 114772 9602
rect 114716 8708 114772 9550
rect 114828 9266 114884 9998
rect 114940 9604 114996 15092
rect 115052 10836 115108 20748
rect 116956 20188 117012 102452
rect 116508 20132 117012 20188
rect 118300 24164 118356 24174
rect 115836 19348 115892 19358
rect 115276 14420 115332 14430
rect 115276 11506 115332 14364
rect 115276 11454 115278 11506
rect 115330 11454 115332 11506
rect 115276 11172 115332 11454
rect 115276 11106 115332 11116
rect 115500 11844 115556 11854
rect 115388 10836 115444 10846
rect 115052 10834 115444 10836
rect 115052 10782 115054 10834
rect 115106 10782 115390 10834
rect 115442 10782 115444 10834
rect 115052 10780 115444 10782
rect 115052 10770 115108 10780
rect 115164 9940 115220 9950
rect 115052 9604 115108 9614
rect 114940 9602 115108 9604
rect 114940 9550 115054 9602
rect 115106 9550 115108 9602
rect 114940 9548 115108 9550
rect 114828 9214 114830 9266
rect 114882 9214 114884 9266
rect 114828 9202 114884 9214
rect 114940 9268 114996 9278
rect 114716 8642 114772 8652
rect 114156 8036 114212 8046
rect 114156 7942 114212 7980
rect 114380 7700 114436 7710
rect 114380 7606 114436 7644
rect 114268 7364 114324 7374
rect 114044 6468 114100 6636
rect 113708 5394 113764 5404
rect 113820 6412 114100 6468
rect 114156 7252 114212 7262
rect 113820 5572 113876 6412
rect 114044 6132 114100 6142
rect 114044 6038 114100 6076
rect 113036 5170 113092 5180
rect 113820 5234 113876 5516
rect 113820 5182 113822 5234
rect 113874 5182 113876 5234
rect 113820 5170 113876 5182
rect 113932 5460 113988 5470
rect 113932 5122 113988 5404
rect 113932 5070 113934 5122
rect 113986 5070 113988 5122
rect 113932 5058 113988 5070
rect 113036 5012 113092 5022
rect 113036 5010 113876 5012
rect 113036 4958 113038 5010
rect 113090 4958 113876 5010
rect 113036 4956 113876 4958
rect 113036 4946 113092 4956
rect 113372 4676 113428 4686
rect 112812 4508 112980 4564
rect 113260 4564 113316 4574
rect 112812 3554 112868 4508
rect 113260 4470 113316 4508
rect 113372 4562 113428 4620
rect 113372 4510 113374 4562
rect 113426 4510 113428 4562
rect 113372 4498 113428 4510
rect 113708 4564 113764 4574
rect 113708 4338 113764 4508
rect 113820 4450 113876 4956
rect 113932 4900 113988 4910
rect 113932 4562 113988 4844
rect 113932 4510 113934 4562
rect 113986 4510 113988 4562
rect 113932 4498 113988 4510
rect 113820 4398 113822 4450
rect 113874 4398 113876 4450
rect 113820 4386 113876 4398
rect 113708 4286 113710 4338
rect 113762 4286 113764 4338
rect 113708 4274 113764 4286
rect 114156 4338 114212 7196
rect 114268 6468 114324 7308
rect 114380 6804 114436 6814
rect 114492 6804 114548 8428
rect 114716 8260 114772 8270
rect 114716 7700 114772 8204
rect 114940 8258 114996 9212
rect 114940 8206 114942 8258
rect 114994 8206 114996 8258
rect 114940 8194 114996 8206
rect 114716 7634 114772 7644
rect 114828 8036 114884 8046
rect 114828 7698 114884 7980
rect 114828 7646 114830 7698
rect 114882 7646 114884 7698
rect 114828 7634 114884 7646
rect 114380 6802 114548 6804
rect 114380 6750 114382 6802
rect 114434 6750 114548 6802
rect 114380 6748 114548 6750
rect 114716 7476 114772 7486
rect 114380 6738 114436 6748
rect 114268 6132 114324 6412
rect 114380 6132 114436 6142
rect 114268 6130 114436 6132
rect 114268 6078 114382 6130
rect 114434 6078 114436 6130
rect 114268 6076 114436 6078
rect 114380 6066 114436 6076
rect 114604 5010 114660 5022
rect 114604 4958 114606 5010
rect 114658 4958 114660 5010
rect 114604 4452 114660 4958
rect 114604 4386 114660 4396
rect 114156 4286 114158 4338
rect 114210 4286 114212 4338
rect 114156 4274 114212 4286
rect 114492 4228 114548 4238
rect 112812 3502 112814 3554
rect 112866 3502 112868 3554
rect 112812 3490 112868 3502
rect 112924 3668 112980 3678
rect 112700 2706 112756 2716
rect 111804 1362 111860 1372
rect 112924 800 112980 3612
rect 114044 3668 114100 3678
rect 114044 3574 114100 3612
rect 113372 3556 113428 3566
rect 113372 3462 113428 3500
rect 114492 1428 114548 4172
rect 114492 1362 114548 1372
rect 114604 3444 114660 3454
rect 114604 800 114660 3388
rect 114716 2212 114772 7420
rect 114828 6466 114884 6478
rect 114828 6414 114830 6466
rect 114882 6414 114884 6466
rect 114828 6356 114884 6414
rect 114828 5124 114884 6300
rect 115052 6244 115108 9548
rect 115164 8260 115220 9884
rect 115164 8194 115220 8204
rect 115164 8034 115220 8046
rect 115164 7982 115166 8034
rect 115218 7982 115220 8034
rect 115164 7252 115220 7982
rect 115164 7186 115220 7196
rect 115052 6178 115108 6188
rect 115164 7028 115220 7038
rect 114828 5058 114884 5068
rect 114940 6020 114996 6030
rect 114940 5348 114996 5964
rect 114940 4562 114996 5292
rect 114940 4510 114942 4562
rect 114994 4510 114996 4562
rect 114940 4498 114996 4510
rect 115164 4228 115220 6972
rect 115276 6018 115332 10780
rect 115388 10770 115444 10780
rect 115500 10050 115556 11788
rect 115500 9998 115502 10050
rect 115554 9998 115556 10050
rect 115500 9828 115556 9998
rect 115388 9772 115556 9828
rect 115612 10724 115668 10734
rect 115388 9154 115444 9772
rect 115388 9102 115390 9154
rect 115442 9102 115444 9154
rect 115388 9090 115444 9102
rect 115500 9602 115556 9614
rect 115500 9550 115502 9602
rect 115554 9550 115556 9602
rect 115500 9380 115556 9550
rect 115500 9044 115556 9324
rect 115500 8978 115556 8988
rect 115612 7924 115668 10668
rect 115836 9268 115892 19292
rect 116396 15876 116452 15886
rect 115948 10498 116004 10510
rect 115948 10446 115950 10498
rect 116002 10446 116004 10498
rect 115948 10164 116004 10446
rect 115948 10098 116004 10108
rect 116060 10388 116116 10398
rect 116060 9940 116116 10332
rect 116396 10052 116452 15820
rect 116060 9938 116340 9940
rect 116060 9886 116062 9938
rect 116114 9886 116340 9938
rect 116060 9884 116340 9886
rect 116060 9874 116116 9884
rect 115836 9202 115892 9212
rect 115948 9380 116004 9390
rect 115724 9154 115780 9166
rect 115724 9102 115726 9154
rect 115778 9102 115780 9154
rect 115724 8372 115780 9102
rect 115724 8306 115780 8316
rect 115836 8932 115892 8942
rect 115500 7868 115668 7924
rect 115724 8036 115780 8046
rect 115388 7476 115444 7486
rect 115388 7382 115444 7420
rect 115500 7028 115556 7868
rect 115500 6962 115556 6972
rect 115612 7474 115668 7486
rect 115612 7422 115614 7474
rect 115666 7422 115668 7474
rect 115500 6804 115556 6814
rect 115612 6804 115668 7422
rect 115724 7476 115780 7980
rect 115836 7698 115892 8876
rect 115948 8036 116004 9324
rect 116284 9156 116340 9884
rect 116060 9154 116340 9156
rect 116060 9102 116286 9154
rect 116338 9102 116340 9154
rect 116060 9100 116340 9102
rect 116060 8260 116116 9100
rect 116284 9090 116340 9100
rect 116396 9156 116452 9996
rect 116396 9090 116452 9100
rect 116060 8128 116116 8204
rect 116508 8148 116564 20132
rect 117180 12068 117236 12078
rect 116732 11172 116788 11182
rect 116732 10834 116788 11116
rect 116732 10782 116734 10834
rect 116786 10782 116788 10834
rect 116620 9716 116676 9726
rect 116620 9266 116676 9660
rect 116620 9214 116622 9266
rect 116674 9214 116676 9266
rect 116620 9202 116676 9214
rect 116732 8708 116788 10782
rect 117180 9826 117236 12012
rect 117404 10836 117460 10846
rect 117292 10500 117348 10510
rect 117292 10406 117348 10444
rect 117180 9774 117182 9826
rect 117234 9774 117236 9826
rect 117180 9762 117236 9774
rect 117068 9716 117124 9726
rect 116732 8642 116788 8652
rect 116844 9714 117124 9716
rect 116844 9662 117070 9714
rect 117122 9662 117124 9714
rect 116844 9660 117124 9662
rect 116508 8082 116564 8092
rect 116732 8148 116788 8158
rect 115948 7980 116116 8036
rect 115836 7646 115838 7698
rect 115890 7646 115892 7698
rect 115836 7634 115892 7646
rect 115948 7588 116004 7598
rect 115948 7494 116004 7532
rect 115724 7410 115780 7420
rect 115500 6802 115668 6804
rect 115500 6750 115502 6802
rect 115554 6750 115668 6802
rect 115500 6748 115668 6750
rect 115836 7252 115892 7262
rect 115500 6738 115556 6748
rect 115724 6578 115780 6590
rect 115724 6526 115726 6578
rect 115778 6526 115780 6578
rect 115276 5966 115278 6018
rect 115330 5966 115332 6018
rect 115276 5122 115332 5966
rect 115276 5070 115278 5122
rect 115330 5070 115332 5122
rect 115276 5058 115332 5070
rect 115612 6018 115668 6030
rect 115612 5966 115614 6018
rect 115666 5966 115668 6018
rect 115500 4898 115556 4910
rect 115500 4846 115502 4898
rect 115554 4846 115556 4898
rect 115500 4676 115556 4846
rect 115612 4900 115668 5966
rect 115724 5124 115780 6526
rect 115724 5058 115780 5068
rect 115612 4834 115668 4844
rect 115724 4676 115780 4686
rect 115500 4620 115724 4676
rect 115724 4562 115780 4620
rect 115724 4510 115726 4562
rect 115778 4510 115780 4562
rect 115724 4498 115780 4510
rect 115164 4162 115220 4172
rect 115500 4338 115556 4350
rect 115500 4286 115502 4338
rect 115554 4286 115556 4338
rect 115500 4228 115556 4286
rect 115500 4162 115556 4172
rect 115724 3556 115780 3566
rect 115836 3556 115892 7196
rect 115948 6692 116004 6702
rect 115948 6578 116004 6636
rect 115948 6526 115950 6578
rect 116002 6526 116004 6578
rect 115948 6514 116004 6526
rect 116060 6578 116116 7980
rect 116060 6526 116062 6578
rect 116114 6526 116116 6578
rect 116060 6514 116116 6526
rect 116172 7924 116228 7934
rect 116060 6132 116116 6142
rect 116172 6132 116228 7868
rect 116396 7362 116452 7374
rect 116396 7310 116398 7362
rect 116450 7310 116452 7362
rect 116284 6468 116340 6478
rect 116284 6374 116340 6412
rect 116060 6130 116228 6132
rect 116060 6078 116062 6130
rect 116114 6078 116228 6130
rect 116060 6076 116228 6078
rect 116060 6066 116116 6076
rect 116396 6020 116452 7310
rect 116396 5954 116452 5964
rect 116620 6692 116676 6702
rect 116508 5796 116564 5806
rect 116396 5794 116564 5796
rect 116396 5742 116510 5794
rect 116562 5742 116564 5794
rect 116396 5740 116564 5742
rect 116060 5348 116116 5358
rect 115948 4898 116004 4910
rect 115948 4846 115950 4898
rect 116002 4846 116004 4898
rect 115948 4788 116004 4846
rect 115948 4722 116004 4732
rect 116060 4564 116116 5292
rect 116060 4338 116116 4508
rect 116172 4452 116228 4462
rect 116172 4358 116228 4396
rect 116060 4286 116062 4338
rect 116114 4286 116116 4338
rect 116060 4274 116116 4286
rect 116396 3892 116452 5740
rect 116508 5730 116564 5740
rect 116508 4340 116564 4350
rect 116620 4340 116676 6636
rect 116508 4338 116676 4340
rect 116508 4286 116510 4338
rect 116562 4286 116676 4338
rect 116508 4284 116676 4286
rect 116732 4338 116788 8092
rect 116844 4562 116900 9660
rect 117068 9650 117124 9660
rect 117292 9716 117348 9754
rect 117292 9650 117348 9660
rect 117404 9492 117460 10780
rect 117068 9436 117460 9492
rect 117740 10498 117796 10510
rect 118188 10500 118244 10576
rect 117740 10446 117742 10498
rect 117794 10446 117796 10498
rect 116956 8260 117012 8270
rect 116956 8166 117012 8204
rect 117068 6466 117124 9436
rect 117180 9156 117236 9166
rect 117180 8932 117236 9100
rect 117516 9156 117572 9166
rect 117516 9062 117572 9100
rect 117180 8876 117572 8932
rect 117404 8708 117460 8718
rect 117292 8596 117348 8606
rect 117068 6414 117070 6466
rect 117122 6414 117124 6466
rect 116956 6356 117012 6366
rect 116956 6130 117012 6300
rect 116956 6078 116958 6130
rect 117010 6078 117012 6130
rect 116956 6066 117012 6078
rect 117068 5908 117124 6414
rect 116844 4510 116846 4562
rect 116898 4510 116900 4562
rect 116844 4498 116900 4510
rect 116956 5852 117124 5908
rect 117180 8372 117236 8382
rect 116732 4286 116734 4338
rect 116786 4286 116788 4338
rect 116508 4274 116564 4284
rect 116732 4274 116788 4286
rect 116956 4116 117012 5852
rect 117068 5348 117124 5358
rect 117068 5010 117124 5292
rect 117068 4958 117070 5010
rect 117122 4958 117124 5010
rect 117068 4946 117124 4958
rect 116956 4050 117012 4060
rect 116396 3826 116452 3836
rect 115724 3554 115892 3556
rect 115724 3502 115726 3554
rect 115778 3502 115892 3554
rect 115724 3500 115892 3502
rect 116284 3668 116340 3678
rect 115724 3490 115780 3500
rect 114716 2146 114772 2156
rect 116284 800 116340 3612
rect 117180 3556 117236 8316
rect 117292 7474 117348 8540
rect 117292 7422 117294 7474
rect 117346 7422 117348 7474
rect 117292 7140 117348 7422
rect 117292 7074 117348 7084
rect 117404 7028 117460 8652
rect 117516 8370 117572 8876
rect 117516 8318 117518 8370
rect 117570 8318 117572 8370
rect 117516 8306 117572 8318
rect 117628 7586 117684 7598
rect 117628 7534 117630 7586
rect 117682 7534 117684 7586
rect 117628 7476 117684 7534
rect 117628 7410 117684 7420
rect 117404 6972 117572 7028
rect 117404 6804 117460 6814
rect 117404 6690 117460 6748
rect 117404 6638 117406 6690
rect 117458 6638 117460 6690
rect 117404 6626 117460 6638
rect 117516 6020 117572 6972
rect 117740 6580 117796 10446
rect 118076 10444 118188 10500
rect 117964 8932 118020 8942
rect 117964 8484 118020 8876
rect 117852 8034 117908 8046
rect 117852 7982 117854 8034
rect 117906 7982 117908 8034
rect 117852 6804 117908 7982
rect 117964 7700 118020 8428
rect 118076 8148 118132 10444
rect 118188 10434 118244 10444
rect 118188 10276 118244 10286
rect 118188 10050 118244 10220
rect 118188 9998 118190 10050
rect 118242 9998 118244 10050
rect 118188 9986 118244 9998
rect 118300 9828 118356 24108
rect 118076 8082 118132 8092
rect 118188 9772 118356 9828
rect 118188 7812 118244 9772
rect 118412 9716 118468 9726
rect 118300 9660 118412 9716
rect 118300 9602 118356 9660
rect 118300 9550 118302 9602
rect 118354 9550 118356 9602
rect 118300 9538 118356 9550
rect 118412 9042 118468 9660
rect 118412 8990 118414 9042
rect 118466 8990 118468 9042
rect 118412 8978 118468 8990
rect 118524 9714 118580 9726
rect 118524 9662 118526 9714
rect 118578 9662 118580 9714
rect 118300 8036 118356 8046
rect 118300 7942 118356 7980
rect 118412 7812 118468 7822
rect 118188 7756 118356 7812
rect 117964 7644 118244 7700
rect 118188 7586 118244 7644
rect 118188 7534 118190 7586
rect 118242 7534 118244 7586
rect 118188 7522 118244 7534
rect 117852 6738 117908 6748
rect 118188 7252 118244 7262
rect 117628 6524 117796 6580
rect 117852 6580 117908 6590
rect 117852 6578 118132 6580
rect 117852 6526 117854 6578
rect 117906 6526 118132 6578
rect 117852 6524 118132 6526
rect 117628 6244 117684 6524
rect 117852 6514 117908 6524
rect 117628 6188 118020 6244
rect 117628 6020 117684 6030
rect 117516 5964 117628 6020
rect 117516 5348 117572 5964
rect 117628 5888 117684 5964
rect 117740 5684 117796 5694
rect 117740 5590 117796 5628
rect 117516 5282 117572 5292
rect 117404 5124 117460 5134
rect 117460 5068 117684 5124
rect 117404 5010 117460 5068
rect 117404 4958 117406 5010
rect 117458 4958 117460 5010
rect 117404 4946 117460 4958
rect 117516 4900 117572 4910
rect 117404 4564 117460 4574
rect 117404 4470 117460 4508
rect 117516 4562 117572 4844
rect 117516 4510 117518 4562
rect 117570 4510 117572 4562
rect 117516 4498 117572 4510
rect 117628 4788 117684 5068
rect 117628 4338 117684 4732
rect 117628 4286 117630 4338
rect 117682 4286 117684 4338
rect 117628 4274 117684 4286
rect 117964 4450 118020 6188
rect 118076 5908 118132 6524
rect 118076 5842 118132 5852
rect 117964 4398 117966 4450
rect 118018 4398 118020 4450
rect 117964 4340 118020 4398
rect 117964 4274 118020 4284
rect 118076 4562 118132 4574
rect 118076 4510 118078 4562
rect 118130 4510 118132 4562
rect 117964 3668 118020 3678
rect 117964 3574 118020 3612
rect 117292 3556 117348 3566
rect 117180 3554 117348 3556
rect 117180 3502 117294 3554
rect 117346 3502 117348 3554
rect 117180 3500 117348 3502
rect 117292 3490 117348 3500
rect 116396 3444 116452 3482
rect 116396 3378 116452 3388
rect 117964 3444 118020 3454
rect 117964 800 118020 3388
rect 118076 3332 118132 4510
rect 118188 4226 118244 7196
rect 118300 5010 118356 7756
rect 118412 7586 118468 7756
rect 118524 7700 118580 9662
rect 118636 9604 118692 9614
rect 118636 9266 118692 9548
rect 118636 9214 118638 9266
rect 118690 9214 118692 9266
rect 118636 9202 118692 9214
rect 118748 8818 118804 8830
rect 118748 8766 118750 8818
rect 118802 8766 118804 8818
rect 118748 8372 118804 8766
rect 118748 8306 118804 8316
rect 118524 7634 118580 7644
rect 118748 8036 118804 8046
rect 118412 7534 118414 7586
rect 118466 7534 118468 7586
rect 118412 7522 118468 7534
rect 118524 7476 118580 7486
rect 118412 5908 118468 5918
rect 118524 5908 118580 7420
rect 118748 7476 118804 7980
rect 118860 8034 118916 8046
rect 118860 7982 118862 8034
rect 118914 7982 118916 8034
rect 118860 7924 118916 7982
rect 118860 7588 118916 7868
rect 118860 7522 118916 7532
rect 118412 5906 118580 5908
rect 118412 5854 118414 5906
rect 118466 5854 118580 5906
rect 118412 5852 118580 5854
rect 118636 7362 118692 7374
rect 118636 7310 118638 7362
rect 118690 7310 118692 7362
rect 118748 7344 118804 7420
rect 118972 7364 119028 116172
rect 120092 11844 120148 116396
rect 120988 116450 121044 116462
rect 120988 116398 120990 116450
rect 121042 116398 121044 116450
rect 120988 115892 121044 116398
rect 123340 116450 123396 116462
rect 123340 116398 123342 116450
rect 123394 116398 123396 116450
rect 122556 116228 122612 116238
rect 122556 116134 122612 116172
rect 123340 116228 123396 116398
rect 123340 116162 123396 116172
rect 125244 116450 125300 116462
rect 127260 116452 127316 116462
rect 125244 116398 125246 116450
rect 125298 116398 125300 116450
rect 121100 115892 121156 115902
rect 120988 115890 121156 115892
rect 120988 115838 121102 115890
rect 121154 115838 121156 115890
rect 120988 115836 121156 115838
rect 121100 115826 121156 115836
rect 125132 115892 125188 115902
rect 125244 115892 125300 116398
rect 125132 115890 125300 115892
rect 125132 115838 125134 115890
rect 125186 115838 125300 115890
rect 125132 115836 125300 115838
rect 126924 116450 127316 116452
rect 126924 116398 127262 116450
rect 127314 116398 127316 116450
rect 126924 116396 127316 116398
rect 126924 115890 126980 116396
rect 127260 116386 127316 116396
rect 129836 116452 129892 116462
rect 126924 115838 126926 115890
rect 126978 115838 126980 115890
rect 125132 115826 125188 115836
rect 120316 115668 120372 115678
rect 120316 115574 120372 115612
rect 121324 115668 121380 115678
rect 121324 115574 121380 115612
rect 124236 115668 124292 115678
rect 124236 115574 124292 115612
rect 124796 115668 124852 115678
rect 124796 115574 124852 115612
rect 125244 115556 125300 115566
rect 120540 27076 120596 27086
rect 120540 15148 120596 27020
rect 120764 26964 120820 26974
rect 120764 20188 120820 26908
rect 124572 24052 124628 24062
rect 123340 22260 123396 22270
rect 120764 20132 120932 20188
rect 120092 11778 120148 11788
rect 120428 15092 120596 15148
rect 119308 11172 119364 11182
rect 119084 11060 119140 11070
rect 119084 10050 119140 11004
rect 119084 9998 119086 10050
rect 119138 9998 119140 10050
rect 119084 9986 119140 9998
rect 119308 10052 119364 11116
rect 120204 10724 120260 10734
rect 119308 9986 119364 9996
rect 119980 10388 120036 10398
rect 119196 9716 119252 9726
rect 119196 9622 119252 9660
rect 119420 9714 119476 9726
rect 119420 9662 119422 9714
rect 119474 9662 119476 9714
rect 119308 9156 119364 9166
rect 119196 8932 119252 8942
rect 119084 8876 119196 8932
rect 119084 8260 119140 8876
rect 119196 8838 119252 8876
rect 119084 8194 119140 8204
rect 119196 8708 119252 8718
rect 118636 5908 118692 7310
rect 118972 7298 119028 7308
rect 118972 7140 119028 7150
rect 118748 6468 118804 6478
rect 118748 6374 118804 6412
rect 118412 5842 118468 5852
rect 118636 5842 118692 5852
rect 118524 5682 118580 5694
rect 118524 5630 118526 5682
rect 118578 5630 118580 5682
rect 118524 5124 118580 5630
rect 118748 5684 118804 5694
rect 118748 5590 118804 5628
rect 118860 5682 118916 5694
rect 118860 5630 118862 5682
rect 118914 5630 118916 5682
rect 118524 5058 118580 5068
rect 118636 5572 118692 5582
rect 118300 4958 118302 5010
rect 118354 4958 118356 5010
rect 118300 4946 118356 4958
rect 118636 5010 118692 5516
rect 118636 4958 118638 5010
rect 118690 4958 118692 5010
rect 118636 4946 118692 4958
rect 118860 4340 118916 5630
rect 118972 5124 119028 7084
rect 119084 6804 119140 6814
rect 119084 6710 119140 6748
rect 118972 5058 119028 5068
rect 119084 5572 119140 5582
rect 118860 4274 118916 4284
rect 118188 4174 118190 4226
rect 118242 4174 118244 4226
rect 118188 4162 118244 4174
rect 118636 4228 118692 4238
rect 118636 4134 118692 4172
rect 118076 3266 118132 3276
rect 119084 800 119140 5516
rect 119196 5122 119252 8652
rect 119308 7140 119364 9100
rect 119420 7588 119476 9662
rect 119868 9602 119924 9614
rect 119868 9550 119870 9602
rect 119922 9550 119924 9602
rect 119644 8932 119700 8942
rect 119532 8930 119700 8932
rect 119532 8878 119646 8930
rect 119698 8878 119700 8930
rect 119532 8876 119700 8878
rect 119532 8818 119588 8876
rect 119644 8866 119700 8876
rect 119532 8766 119534 8818
rect 119586 8766 119588 8818
rect 119532 8146 119588 8766
rect 119868 8708 119924 9550
rect 119868 8642 119924 8652
rect 119980 8596 120036 10332
rect 120204 10388 120260 10668
rect 120204 10322 120260 10332
rect 120316 9268 120372 9278
rect 120092 8930 120148 8942
rect 120092 8878 120094 8930
rect 120146 8878 120148 8930
rect 120092 8818 120148 8878
rect 120092 8766 120094 8818
rect 120146 8766 120148 8818
rect 120092 8754 120148 8766
rect 119980 8540 120148 8596
rect 119980 8372 120036 8382
rect 119644 8260 119700 8270
rect 119644 8166 119700 8204
rect 119756 8258 119812 8270
rect 119756 8206 119758 8258
rect 119810 8206 119812 8258
rect 119532 8094 119534 8146
rect 119586 8094 119588 8146
rect 119532 7812 119588 8094
rect 119756 8036 119812 8206
rect 119756 7970 119812 7980
rect 119588 7756 119700 7812
rect 119532 7746 119588 7756
rect 119644 7588 119700 7756
rect 119420 7532 119588 7588
rect 119420 7364 119476 7374
rect 119420 7270 119476 7308
rect 119308 7084 119476 7140
rect 119308 6916 119364 6926
rect 119308 6690 119364 6860
rect 119308 6638 119310 6690
rect 119362 6638 119364 6690
rect 119308 6626 119364 6638
rect 119420 6356 119476 7084
rect 119532 7028 119588 7532
rect 119644 7474 119700 7532
rect 119644 7422 119646 7474
rect 119698 7422 119700 7474
rect 119644 7410 119700 7422
rect 119532 6962 119588 6972
rect 119868 6916 119924 6926
rect 119196 5070 119198 5122
rect 119250 5070 119252 5122
rect 119196 2884 119252 5070
rect 119308 6300 119476 6356
rect 119756 6804 119812 6814
rect 119308 3556 119364 6300
rect 119756 5906 119812 6748
rect 119868 6356 119924 6860
rect 119868 6290 119924 6300
rect 119756 5854 119758 5906
rect 119810 5854 119812 5906
rect 119756 5842 119812 5854
rect 119868 5908 119924 5918
rect 119868 5814 119924 5852
rect 119420 5682 119476 5694
rect 119420 5630 119422 5682
rect 119474 5630 119476 5682
rect 119420 5348 119476 5630
rect 119532 5684 119588 5694
rect 119532 5590 119588 5628
rect 119644 5348 119700 5358
rect 119420 5346 119700 5348
rect 119420 5294 119646 5346
rect 119698 5294 119700 5346
rect 119420 5292 119700 5294
rect 119644 5282 119700 5292
rect 119868 5236 119924 5246
rect 119868 5142 119924 5180
rect 119980 5234 120036 8316
rect 120092 6916 120148 8540
rect 120092 6850 120148 6860
rect 120204 8034 120260 8046
rect 120204 7982 120206 8034
rect 120258 7982 120260 8034
rect 120204 6804 120260 7982
rect 120316 7812 120372 9212
rect 120428 8036 120484 15092
rect 120876 9268 120932 20132
rect 123228 17556 123284 17566
rect 120988 9268 121044 9278
rect 120932 9266 121044 9268
rect 120932 9214 120990 9266
rect 121042 9214 121044 9266
rect 120932 9212 121044 9214
rect 120876 9202 120932 9212
rect 120988 9202 121044 9212
rect 121884 9268 121940 9278
rect 121884 9174 121940 9212
rect 120988 9044 121044 9054
rect 120988 8596 121044 8988
rect 121548 9044 121604 9054
rect 121548 8950 121604 8988
rect 120428 7970 120484 7980
rect 120540 8540 121044 8596
rect 120316 7756 120484 7812
rect 120316 7364 120372 7374
rect 120316 7270 120372 7308
rect 120428 7140 120484 7756
rect 120204 6672 120260 6748
rect 120316 7084 120484 7140
rect 120316 6580 120372 7084
rect 120204 6524 120372 6580
rect 120428 6690 120484 6702
rect 120428 6638 120430 6690
rect 120482 6638 120484 6690
rect 119980 5182 119982 5234
rect 120034 5182 120036 5234
rect 119980 5170 120036 5182
rect 120092 6468 120148 6478
rect 119756 5124 119812 5134
rect 119420 5010 119476 5022
rect 119420 4958 119422 5010
rect 119474 4958 119476 5010
rect 119420 4900 119476 4958
rect 119476 4844 119700 4900
rect 119420 4834 119476 4844
rect 119420 4452 119476 4462
rect 119420 4358 119476 4396
rect 119644 4450 119700 4844
rect 119756 4562 119812 5068
rect 120092 5122 120148 6412
rect 120092 5070 120094 5122
rect 120146 5070 120148 5122
rect 120092 5058 120148 5070
rect 119756 4510 119758 4562
rect 119810 4510 119812 4562
rect 119756 4498 119812 4510
rect 119644 4398 119646 4450
rect 119698 4398 119700 4450
rect 119644 3892 119700 4398
rect 120204 4452 120260 6524
rect 120428 6356 120484 6638
rect 120428 6290 120484 6300
rect 120204 4386 120260 4396
rect 120316 4452 120372 4462
rect 120540 4452 120596 8540
rect 120988 8372 121044 8382
rect 120652 8260 120708 8270
rect 120652 8166 120708 8204
rect 120764 8036 120820 8046
rect 120652 6692 120708 6702
rect 120652 6356 120708 6636
rect 120652 6290 120708 6300
rect 120764 5010 120820 7980
rect 120988 7698 121044 8316
rect 121212 8148 121268 8158
rect 120988 7646 120990 7698
rect 121042 7646 121044 7698
rect 120988 7634 121044 7646
rect 121100 8034 121156 8046
rect 121100 7982 121102 8034
rect 121154 7982 121156 8034
rect 121100 7140 121156 7982
rect 121100 7074 121156 7084
rect 121100 6578 121156 6590
rect 121100 6526 121102 6578
rect 121154 6526 121156 6578
rect 121100 6468 121156 6526
rect 120876 6412 121156 6468
rect 120876 5124 120932 6412
rect 121212 6244 121268 8092
rect 121548 8036 121604 8046
rect 121996 8036 122052 8046
rect 121548 8034 121716 8036
rect 121548 7982 121550 8034
rect 121602 7982 121716 8034
rect 121548 7980 121716 7982
rect 121548 7970 121604 7980
rect 121436 7588 121492 7598
rect 121436 7494 121492 7532
rect 120876 5058 120932 5068
rect 120988 6188 121268 6244
rect 121324 7364 121380 7374
rect 120764 4958 120766 5010
rect 120818 4958 120820 5010
rect 120764 4946 120820 4958
rect 120876 4898 120932 4910
rect 120876 4846 120878 4898
rect 120930 4846 120932 4898
rect 120876 4564 120932 4846
rect 120876 4498 120932 4508
rect 120316 4450 120596 4452
rect 120316 4398 120318 4450
rect 120370 4398 120596 4450
rect 120316 4396 120596 4398
rect 120316 4386 120372 4396
rect 119868 4340 119924 4350
rect 119868 4246 119924 4284
rect 119644 3826 119700 3836
rect 120092 4226 120148 4238
rect 120092 4174 120094 4226
rect 120146 4174 120148 4226
rect 119420 3556 119476 3566
rect 119308 3554 119476 3556
rect 119308 3502 119422 3554
rect 119474 3502 119476 3554
rect 119308 3500 119476 3502
rect 119420 3490 119476 3500
rect 119196 2818 119252 2828
rect 119644 3332 119700 3342
rect 119644 800 119700 3276
rect 120092 3108 120148 4174
rect 120092 3042 120148 3052
rect 120204 3780 120260 3790
rect 120204 800 120260 3724
rect 120764 3668 120820 3678
rect 120316 3444 120372 3482
rect 120316 3378 120372 3388
rect 120764 800 120820 3612
rect 120988 3444 121044 6188
rect 121212 6018 121268 6030
rect 121212 5966 121214 6018
rect 121266 5966 121268 6018
rect 121100 5796 121156 5806
rect 121100 5702 121156 5740
rect 121212 5348 121268 5966
rect 121100 5292 121268 5348
rect 121100 4900 121156 5292
rect 121100 4834 121156 4844
rect 121212 5122 121268 5134
rect 121212 5070 121214 5122
rect 121266 5070 121268 5122
rect 121212 4676 121268 5070
rect 121324 5010 121380 7308
rect 121548 6466 121604 6478
rect 121548 6414 121550 6466
rect 121602 6414 121604 6466
rect 121436 5796 121492 5806
rect 121436 5702 121492 5740
rect 121324 4958 121326 5010
rect 121378 4958 121380 5010
rect 121324 4946 121380 4958
rect 121212 4610 121268 4620
rect 121436 4676 121492 4686
rect 121324 4564 121380 4574
rect 121324 4470 121380 4508
rect 121212 4340 121268 4350
rect 121212 4246 121268 4284
rect 121436 4338 121492 4620
rect 121548 4452 121604 6414
rect 121660 5572 121716 7980
rect 121996 7942 122052 7980
rect 122556 8034 122612 8046
rect 122556 7982 122558 8034
rect 122610 7982 122612 8034
rect 121884 7924 121940 7934
rect 121660 5506 121716 5516
rect 121772 7028 121828 7038
rect 121660 5348 121716 5358
rect 121660 5234 121716 5292
rect 121660 5182 121662 5234
rect 121714 5182 121716 5234
rect 121660 5170 121716 5182
rect 121772 5234 121828 6972
rect 121884 5460 121940 7868
rect 122220 7812 122276 7822
rect 121996 7364 122052 7374
rect 121996 6916 122052 7308
rect 121996 6850 122052 6860
rect 121996 6468 122052 6478
rect 121996 6020 122052 6412
rect 121996 5954 122052 5964
rect 121996 5796 122052 5806
rect 121996 5702 122052 5740
rect 122108 5794 122164 5806
rect 122108 5742 122110 5794
rect 122162 5742 122164 5794
rect 122108 5460 122164 5742
rect 121884 5404 122052 5460
rect 121772 5182 121774 5234
rect 121826 5182 121828 5234
rect 121772 5170 121828 5182
rect 121884 5236 121940 5246
rect 121884 5142 121940 5180
rect 121772 5012 121828 5022
rect 121548 4386 121604 4396
rect 121660 4564 121716 4574
rect 121436 4286 121438 4338
rect 121490 4286 121492 4338
rect 121436 4274 121492 4286
rect 121548 4116 121604 4126
rect 121436 3892 121492 3902
rect 121212 3556 121268 3566
rect 121212 3462 121268 3500
rect 121436 3554 121492 3836
rect 121436 3502 121438 3554
rect 121490 3502 121492 3554
rect 121436 3490 121492 3502
rect 120988 3378 121044 3388
rect 121548 2436 121604 4060
rect 121660 3554 121716 4508
rect 121772 4450 121828 4956
rect 121772 4398 121774 4450
rect 121826 4398 121828 4450
rect 121772 4386 121828 4398
rect 121996 4116 122052 5404
rect 122108 5394 122164 5404
rect 122108 5012 122164 5022
rect 122108 4338 122164 4956
rect 122220 4562 122276 7756
rect 122556 7700 122612 7982
rect 123004 8034 123060 8046
rect 123004 7982 123006 8034
rect 123058 7982 123060 8034
rect 123004 7924 123060 7982
rect 122332 7644 122612 7700
rect 122780 7868 123060 7924
rect 122332 6132 122388 7644
rect 122444 7476 122500 7486
rect 122780 7476 122836 7868
rect 123228 7700 123284 17500
rect 123228 7568 123284 7644
rect 122444 7362 122500 7420
rect 122444 7310 122446 7362
rect 122498 7310 122500 7362
rect 122444 7252 122500 7310
rect 122444 7186 122500 7196
rect 122668 7420 122836 7476
rect 122444 6692 122500 6702
rect 122444 6598 122500 6636
rect 122332 6066 122388 6076
rect 122332 5906 122388 5918
rect 122332 5854 122334 5906
rect 122386 5854 122388 5906
rect 122332 4676 122388 5854
rect 122668 5908 122724 7420
rect 122892 7364 122948 7374
rect 123340 7364 123396 22204
rect 122892 7362 123060 7364
rect 122892 7310 122894 7362
rect 122946 7310 123060 7362
rect 122892 7308 123060 7310
rect 122892 7298 122948 7308
rect 122892 6804 122948 6814
rect 122780 6802 122948 6804
rect 122780 6750 122894 6802
rect 122946 6750 122948 6802
rect 122780 6748 122948 6750
rect 122780 6692 122836 6748
rect 122892 6738 122948 6748
rect 122780 6626 122836 6636
rect 123004 6580 123060 7308
rect 122892 6524 123060 6580
rect 123116 7308 123396 7364
rect 123452 8932 123508 8942
rect 123452 8370 123508 8876
rect 124124 8820 124180 8830
rect 123452 8318 123454 8370
rect 123506 8318 123508 8370
rect 122668 5348 122724 5852
rect 122668 5282 122724 5292
rect 122780 6468 122836 6478
rect 122444 4900 122500 4910
rect 122444 4898 122612 4900
rect 122444 4846 122446 4898
rect 122498 4846 122612 4898
rect 122444 4844 122612 4846
rect 122444 4834 122500 4844
rect 122556 4788 122612 4844
rect 122556 4732 122724 4788
rect 122332 4620 122612 4676
rect 122220 4510 122222 4562
rect 122274 4510 122276 4562
rect 122220 4498 122276 4510
rect 122108 4286 122110 4338
rect 122162 4286 122164 4338
rect 122108 4274 122164 4286
rect 122332 4340 122388 4350
rect 122332 4246 122388 4284
rect 121772 4060 122052 4116
rect 122220 4228 122276 4238
rect 121772 3666 121828 4060
rect 121772 3614 121774 3666
rect 121826 3614 121828 3666
rect 121772 3602 121828 3614
rect 121884 3668 121940 3678
rect 121660 3502 121662 3554
rect 121714 3502 121716 3554
rect 121660 3490 121716 3502
rect 121772 3444 121828 3482
rect 121772 3378 121828 3388
rect 121324 2380 121604 2436
rect 121324 800 121380 2380
rect 121884 800 121940 3612
rect 122220 3108 122276 4172
rect 122444 3332 122500 3342
rect 122444 3238 122500 3276
rect 122556 3220 122612 4620
rect 122668 4116 122724 4732
rect 122780 4562 122836 6412
rect 122892 5572 122948 6524
rect 123116 6468 123172 7308
rect 123452 6804 123508 8318
rect 123900 8484 123956 8494
rect 123788 8036 123844 8046
rect 123452 6738 123508 6748
rect 123564 8034 123844 8036
rect 123564 7982 123790 8034
rect 123842 7982 123844 8034
rect 123564 7980 123844 7982
rect 123452 6468 123508 6478
rect 122892 5124 122948 5516
rect 123004 6412 123172 6468
rect 123228 6466 123508 6468
rect 123228 6414 123454 6466
rect 123506 6414 123508 6466
rect 123228 6412 123508 6414
rect 123004 5346 123060 6412
rect 123004 5294 123006 5346
rect 123058 5294 123060 5346
rect 123004 5282 123060 5294
rect 123116 6018 123172 6030
rect 123116 5966 123118 6018
rect 123170 5966 123172 6018
rect 122892 5058 122948 5068
rect 122780 4510 122782 4562
rect 122834 4510 122836 4562
rect 122780 4498 122836 4510
rect 122668 4050 122724 4060
rect 122556 3154 122612 3164
rect 122220 3052 122500 3108
rect 122444 800 122500 3052
rect 123116 1540 123172 5966
rect 123004 1484 123172 1540
rect 123228 4004 123284 6412
rect 123452 6402 123508 6412
rect 123340 6132 123396 6142
rect 123340 5124 123396 6076
rect 123452 5348 123508 5358
rect 123452 5254 123508 5292
rect 123340 5068 123508 5124
rect 123004 800 123060 1484
rect 123228 1316 123284 3948
rect 123340 4900 123396 4910
rect 123340 3330 123396 4844
rect 123452 4562 123508 5068
rect 123564 4676 123620 7980
rect 123788 7970 123844 7980
rect 123788 7362 123844 7374
rect 123788 7310 123790 7362
rect 123842 7310 123844 7362
rect 123788 6244 123844 7310
rect 123900 6690 123956 8428
rect 123900 6638 123902 6690
rect 123954 6638 123956 6690
rect 123900 6468 123956 6638
rect 123900 6402 123956 6412
rect 123844 6188 123956 6244
rect 123788 6178 123844 6188
rect 123788 6020 123844 6030
rect 123788 5926 123844 5964
rect 123788 5684 123844 5694
rect 123676 5124 123732 5134
rect 123676 5030 123732 5068
rect 123564 4610 123620 4620
rect 123452 4510 123454 4562
rect 123506 4510 123508 4562
rect 123452 4498 123508 4510
rect 123676 4564 123732 4574
rect 123788 4564 123844 5628
rect 123900 5346 123956 6188
rect 124124 5908 124180 8764
rect 124236 8708 124292 8718
rect 124236 8148 124292 8652
rect 124236 7698 124292 8092
rect 124236 7646 124238 7698
rect 124290 7646 124292 7698
rect 124236 7634 124292 7646
rect 124348 8034 124404 8046
rect 124348 7982 124350 8034
rect 124402 7982 124404 8034
rect 124236 6466 124292 6478
rect 124236 6414 124238 6466
rect 124290 6414 124292 6466
rect 124236 6356 124292 6414
rect 124236 6290 124292 6300
rect 124124 5906 124292 5908
rect 124124 5854 124126 5906
rect 124178 5854 124292 5906
rect 124124 5852 124292 5854
rect 124124 5842 124180 5852
rect 123900 5294 123902 5346
rect 123954 5294 123956 5346
rect 123900 5282 123956 5294
rect 124012 5794 124068 5806
rect 124012 5742 124014 5794
rect 124066 5742 124068 5794
rect 123676 4562 123844 4564
rect 123676 4510 123678 4562
rect 123730 4510 123844 4562
rect 123676 4508 123844 4510
rect 123900 4676 123956 4686
rect 123676 4498 123732 4508
rect 123564 4226 123620 4238
rect 123900 4228 123956 4620
rect 124012 4338 124068 5742
rect 124012 4286 124014 4338
rect 124066 4286 124068 4338
rect 124012 4274 124068 4286
rect 124124 5010 124180 5022
rect 124124 4958 124126 5010
rect 124178 4958 124180 5010
rect 123564 4174 123566 4226
rect 123618 4174 123620 4226
rect 123564 4116 123620 4174
rect 123564 4050 123620 4060
rect 123676 4172 123956 4228
rect 123676 3892 123732 4172
rect 124124 4116 124180 4958
rect 124236 5012 124292 5852
rect 124236 4946 124292 4956
rect 124124 4050 124180 4060
rect 123676 3554 123732 3836
rect 123676 3502 123678 3554
rect 123730 3502 123732 3554
rect 123676 3490 123732 3502
rect 124124 3892 124180 3902
rect 123340 3278 123342 3330
rect 123394 3278 123396 3330
rect 123340 3266 123396 3278
rect 123564 3444 123620 3454
rect 123228 1250 123284 1260
rect 123564 800 123620 3388
rect 124124 800 124180 3836
rect 124348 3556 124404 7982
rect 124460 7250 124516 7262
rect 124460 7198 124462 7250
rect 124514 7198 124516 7250
rect 124460 5348 124516 7198
rect 124460 5282 124516 5292
rect 124572 4562 124628 23996
rect 125244 9940 125300 115500
rect 126924 115556 126980 115838
rect 129836 115890 129892 116396
rect 131180 116452 131236 116462
rect 131180 116358 131236 116396
rect 129836 115838 129838 115890
rect 129890 115838 129892 115890
rect 129836 115826 129892 115838
rect 131516 115780 131572 119200
rect 134652 117010 134708 119200
rect 134652 116958 134654 117010
rect 134706 116958 134708 117010
rect 134652 116946 134708 116958
rect 135772 117010 135828 117022
rect 135772 116958 135774 117010
rect 135826 116958 135828 117010
rect 131852 116564 131908 116574
rect 131852 116470 131908 116508
rect 135772 116562 135828 116958
rect 136220 117010 136276 119200
rect 136220 116958 136222 117010
rect 136274 116958 136276 117010
rect 136220 116946 136276 116958
rect 137564 117010 137620 117022
rect 137564 116958 137566 117010
rect 137618 116958 137620 117010
rect 135772 116510 135774 116562
rect 135826 116510 135828 116562
rect 135772 116498 135828 116510
rect 137564 116562 137620 116958
rect 139356 116676 139412 119200
rect 139356 116610 139412 116620
rect 140252 116676 140308 116686
rect 137564 116510 137566 116562
rect 137618 116510 137620 116562
rect 137564 116498 137620 116510
rect 140252 116562 140308 116620
rect 140252 116510 140254 116562
rect 140306 116510 140308 116562
rect 140252 116498 140308 116510
rect 135100 116452 135156 116462
rect 134652 116450 135156 116452
rect 134652 116398 135102 116450
rect 135154 116398 135156 116450
rect 134652 116396 135156 116398
rect 134652 115890 134708 116396
rect 135100 116386 135156 116396
rect 136892 116450 136948 116462
rect 139580 116452 139636 116462
rect 136892 116398 136894 116450
rect 136946 116398 136948 116450
rect 134652 115838 134654 115890
rect 134706 115838 134708 115890
rect 134652 115826 134708 115838
rect 131516 115714 131572 115724
rect 132636 115780 132692 115790
rect 132636 115686 132692 115724
rect 128940 115668 128996 115678
rect 128940 115574 128996 115612
rect 129612 115668 129668 115678
rect 129612 115574 129668 115612
rect 131740 115666 131796 115678
rect 131740 115614 131742 115666
rect 131794 115614 131796 115666
rect 126924 115490 126980 115500
rect 131292 115556 131348 115566
rect 131740 115556 131796 115614
rect 133756 115668 133812 115678
rect 133756 115574 133812 115612
rect 134316 115668 134372 115678
rect 134316 115574 134372 115612
rect 131292 115554 131796 115556
rect 131292 115502 131294 115554
rect 131346 115502 131796 115554
rect 131292 115500 131796 115502
rect 131292 115490 131348 115500
rect 127356 115276 127620 115286
rect 127412 115220 127460 115276
rect 127516 115220 127564 115276
rect 127356 115210 127620 115220
rect 127356 113708 127620 113718
rect 127412 113652 127460 113708
rect 127516 113652 127564 113708
rect 127356 113642 127620 113652
rect 127356 112140 127620 112150
rect 127412 112084 127460 112140
rect 127516 112084 127564 112140
rect 127356 112074 127620 112084
rect 127356 110572 127620 110582
rect 127412 110516 127460 110572
rect 127516 110516 127564 110572
rect 127356 110506 127620 110516
rect 127356 109004 127620 109014
rect 127412 108948 127460 109004
rect 127516 108948 127564 109004
rect 127356 108938 127620 108948
rect 127356 107436 127620 107446
rect 127412 107380 127460 107436
rect 127516 107380 127564 107436
rect 127356 107370 127620 107380
rect 127356 105868 127620 105878
rect 127412 105812 127460 105868
rect 127516 105812 127564 105868
rect 127356 105802 127620 105812
rect 127356 104300 127620 104310
rect 127412 104244 127460 104300
rect 127516 104244 127564 104300
rect 127356 104234 127620 104244
rect 127356 102732 127620 102742
rect 127412 102676 127460 102732
rect 127516 102676 127564 102732
rect 127356 102666 127620 102676
rect 127356 101164 127620 101174
rect 127412 101108 127460 101164
rect 127516 101108 127564 101164
rect 127356 101098 127620 101108
rect 127356 99596 127620 99606
rect 127412 99540 127460 99596
rect 127516 99540 127564 99596
rect 127356 99530 127620 99540
rect 127356 98028 127620 98038
rect 127412 97972 127460 98028
rect 127516 97972 127564 98028
rect 127356 97962 127620 97972
rect 127356 96460 127620 96470
rect 127412 96404 127460 96460
rect 127516 96404 127564 96460
rect 127356 96394 127620 96404
rect 127356 94892 127620 94902
rect 127412 94836 127460 94892
rect 127516 94836 127564 94892
rect 127356 94826 127620 94836
rect 127356 93324 127620 93334
rect 127412 93268 127460 93324
rect 127516 93268 127564 93324
rect 127356 93258 127620 93268
rect 127356 91756 127620 91766
rect 127412 91700 127460 91756
rect 127516 91700 127564 91756
rect 127356 91690 127620 91700
rect 127356 90188 127620 90198
rect 127412 90132 127460 90188
rect 127516 90132 127564 90188
rect 127356 90122 127620 90132
rect 127356 88620 127620 88630
rect 127412 88564 127460 88620
rect 127516 88564 127564 88620
rect 127356 88554 127620 88564
rect 127356 87052 127620 87062
rect 127412 86996 127460 87052
rect 127516 86996 127564 87052
rect 127356 86986 127620 86996
rect 127356 85484 127620 85494
rect 127412 85428 127460 85484
rect 127516 85428 127564 85484
rect 127356 85418 127620 85428
rect 127356 83916 127620 83926
rect 127412 83860 127460 83916
rect 127516 83860 127564 83916
rect 127356 83850 127620 83860
rect 127356 82348 127620 82358
rect 127412 82292 127460 82348
rect 127516 82292 127564 82348
rect 127356 82282 127620 82292
rect 127356 80780 127620 80790
rect 127412 80724 127460 80780
rect 127516 80724 127564 80780
rect 127356 80714 127620 80724
rect 127356 79212 127620 79222
rect 127412 79156 127460 79212
rect 127516 79156 127564 79212
rect 127356 79146 127620 79156
rect 127356 77644 127620 77654
rect 127412 77588 127460 77644
rect 127516 77588 127564 77644
rect 127356 77578 127620 77588
rect 127356 76076 127620 76086
rect 127412 76020 127460 76076
rect 127516 76020 127564 76076
rect 127356 76010 127620 76020
rect 127356 74508 127620 74518
rect 127412 74452 127460 74508
rect 127516 74452 127564 74508
rect 127356 74442 127620 74452
rect 127356 72940 127620 72950
rect 127412 72884 127460 72940
rect 127516 72884 127564 72940
rect 127356 72874 127620 72884
rect 127356 71372 127620 71382
rect 127412 71316 127460 71372
rect 127516 71316 127564 71372
rect 127356 71306 127620 71316
rect 127356 69804 127620 69814
rect 127412 69748 127460 69804
rect 127516 69748 127564 69804
rect 127356 69738 127620 69748
rect 127356 68236 127620 68246
rect 127412 68180 127460 68236
rect 127516 68180 127564 68236
rect 127356 68170 127620 68180
rect 127356 66668 127620 66678
rect 127412 66612 127460 66668
rect 127516 66612 127564 66668
rect 127356 66602 127620 66612
rect 127356 65100 127620 65110
rect 127412 65044 127460 65100
rect 127516 65044 127564 65100
rect 127356 65034 127620 65044
rect 127356 63532 127620 63542
rect 127412 63476 127460 63532
rect 127516 63476 127564 63532
rect 127356 63466 127620 63476
rect 127356 61964 127620 61974
rect 127412 61908 127460 61964
rect 127516 61908 127564 61964
rect 127356 61898 127620 61908
rect 127356 60396 127620 60406
rect 127412 60340 127460 60396
rect 127516 60340 127564 60396
rect 127356 60330 127620 60340
rect 127356 58828 127620 58838
rect 127412 58772 127460 58828
rect 127516 58772 127564 58828
rect 127356 58762 127620 58772
rect 127356 57260 127620 57270
rect 127412 57204 127460 57260
rect 127516 57204 127564 57260
rect 127356 57194 127620 57204
rect 127356 55692 127620 55702
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127356 55626 127620 55636
rect 127356 54124 127620 54134
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127356 54058 127620 54068
rect 127356 52556 127620 52566
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127356 52490 127620 52500
rect 127356 50988 127620 50998
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127356 50922 127620 50932
rect 127356 49420 127620 49430
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127356 49354 127620 49364
rect 127356 47852 127620 47862
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127356 47786 127620 47796
rect 127356 46284 127620 46294
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127356 46218 127620 46228
rect 127356 44716 127620 44726
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127356 44650 127620 44660
rect 127356 43148 127620 43158
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127356 43082 127620 43092
rect 127356 41580 127620 41590
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127356 41514 127620 41524
rect 127356 40012 127620 40022
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127356 39946 127620 39956
rect 127356 38444 127620 38454
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127356 38378 127620 38388
rect 127356 36876 127620 36886
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127356 36810 127620 36820
rect 127356 35308 127620 35318
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127356 35242 127620 35252
rect 127356 33740 127620 33750
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127356 33674 127620 33684
rect 127356 32172 127620 32182
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127356 32106 127620 32116
rect 127356 30604 127620 30614
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127356 30538 127620 30548
rect 127356 29036 127620 29046
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127356 28970 127620 28980
rect 126364 28644 126420 28654
rect 125244 9874 125300 9884
rect 125692 19236 125748 19246
rect 124684 7362 124740 7374
rect 125020 7364 125076 7374
rect 125468 7364 125524 7374
rect 124684 7310 124686 7362
rect 124738 7310 124740 7362
rect 124684 7250 124740 7310
rect 124684 7198 124686 7250
rect 124738 7198 124740 7250
rect 124684 7186 124740 7198
rect 124796 7362 125076 7364
rect 124796 7310 125022 7362
rect 125074 7310 125076 7362
rect 124796 7308 125076 7310
rect 124796 6356 124852 7308
rect 125020 7298 125076 7308
rect 125244 7362 125524 7364
rect 125244 7310 125470 7362
rect 125522 7310 125524 7362
rect 125244 7308 125524 7310
rect 124908 6468 124964 6478
rect 124908 6466 125188 6468
rect 124908 6414 124910 6466
rect 124962 6414 125188 6466
rect 124908 6412 125188 6414
rect 124908 6402 124964 6412
rect 124796 6290 124852 6300
rect 124908 6020 124964 6030
rect 124572 4510 124574 4562
rect 124626 4510 124628 4562
rect 124572 4498 124628 4510
rect 124684 6018 124964 6020
rect 124684 5966 124910 6018
rect 124962 5966 124964 6018
rect 124684 5964 124964 5966
rect 124460 3556 124516 3566
rect 124404 3554 124516 3556
rect 124404 3502 124462 3554
rect 124514 3502 124516 3554
rect 124404 3500 124516 3502
rect 124348 3424 124404 3500
rect 124460 3490 124516 3500
rect 124236 3332 124292 3342
rect 124236 3238 124292 3276
rect 124684 800 124740 5964
rect 124908 5954 124964 5964
rect 125020 5796 125076 5806
rect 125020 5236 125076 5740
rect 124908 5124 124964 5134
rect 124908 5030 124964 5068
rect 124796 4338 124852 4350
rect 124796 4286 124798 4338
rect 124850 4286 124852 4338
rect 124796 4228 124852 4286
rect 124796 4162 124852 4172
rect 125020 3388 125076 5180
rect 125132 5012 125188 6412
rect 125132 4116 125188 4956
rect 125244 4676 125300 7308
rect 125468 7298 125524 7308
rect 125692 6692 125748 19180
rect 126140 7362 126196 7374
rect 126140 7310 126142 7362
rect 126194 7310 126196 7362
rect 125692 6626 125748 6636
rect 125916 6692 125972 6702
rect 125356 6466 125412 6478
rect 125804 6468 125860 6478
rect 125356 6414 125358 6466
rect 125410 6414 125412 6466
rect 125356 6020 125412 6414
rect 125692 6466 125860 6468
rect 125692 6414 125806 6466
rect 125858 6414 125860 6466
rect 125692 6412 125860 6414
rect 125412 5964 125524 6020
rect 125356 5954 125412 5964
rect 125356 5124 125412 5134
rect 125356 5030 125412 5068
rect 125244 4620 125412 4676
rect 125132 4050 125188 4060
rect 125356 3668 125412 4620
rect 125468 4226 125524 5964
rect 125580 5796 125636 5806
rect 125580 5702 125636 5740
rect 125580 5460 125636 5470
rect 125580 5346 125636 5404
rect 125580 5294 125582 5346
rect 125634 5294 125636 5346
rect 125580 5282 125636 5294
rect 125468 4174 125470 4226
rect 125522 4174 125524 4226
rect 125468 4162 125524 4174
rect 125580 4450 125636 4462
rect 125580 4398 125582 4450
rect 125634 4398 125636 4450
rect 124908 3332 125076 3388
rect 125244 3556 125300 3566
rect 124908 2996 124964 3332
rect 125132 3330 125188 3342
rect 125132 3278 125134 3330
rect 125186 3278 125188 3330
rect 125132 3220 125188 3278
rect 125132 3154 125188 3164
rect 124908 2930 124964 2940
rect 125244 800 125300 3500
rect 125356 3554 125412 3612
rect 125356 3502 125358 3554
rect 125410 3502 125412 3554
rect 125356 3490 125412 3502
rect 125580 3332 125636 4398
rect 125692 4228 125748 6412
rect 125804 6402 125860 6412
rect 125804 6020 125860 6030
rect 125804 5572 125860 5964
rect 125804 5346 125860 5516
rect 125916 5460 125972 6636
rect 126028 5794 126084 5806
rect 126028 5742 126030 5794
rect 126082 5742 126084 5794
rect 126028 5682 126084 5742
rect 126028 5630 126030 5682
rect 126082 5630 126084 5682
rect 126028 5618 126084 5630
rect 125916 5394 125972 5404
rect 125804 5294 125806 5346
rect 125858 5294 125860 5346
rect 125804 5124 125860 5294
rect 126028 5236 126084 5246
rect 126028 5142 126084 5180
rect 125804 5068 125972 5124
rect 125916 5012 125972 5068
rect 125916 4956 126084 5012
rect 125804 4452 125860 4462
rect 125804 4358 125860 4396
rect 125692 4162 125748 4172
rect 125580 3266 125636 3276
rect 125804 3668 125860 3678
rect 126028 3668 126084 4956
rect 126140 3892 126196 7310
rect 126140 3826 126196 3836
rect 126252 5682 126308 5694
rect 126252 5630 126254 5682
rect 126306 5630 126308 5682
rect 126252 4340 126308 5630
rect 126364 4562 126420 28588
rect 127356 27468 127620 27478
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127356 27402 127620 27412
rect 127356 25900 127620 25910
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127356 25834 127620 25844
rect 127356 24332 127620 24342
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127356 24266 127620 24276
rect 127356 22764 127620 22774
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127356 22698 127620 22708
rect 130396 22148 130452 22158
rect 127356 21196 127620 21206
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127356 21130 127620 21140
rect 127148 20692 127204 20702
rect 126476 7364 126532 7374
rect 126476 7362 126644 7364
rect 126476 7310 126478 7362
rect 126530 7310 126644 7362
rect 126476 7308 126644 7310
rect 126476 7298 126532 7308
rect 126476 6466 126532 6478
rect 126476 6414 126478 6466
rect 126530 6414 126532 6466
rect 126476 6020 126532 6414
rect 126476 5954 126532 5964
rect 126476 5794 126532 5806
rect 126476 5742 126478 5794
rect 126530 5742 126532 5794
rect 126476 5682 126532 5742
rect 126476 5630 126478 5682
rect 126530 5630 126532 5682
rect 126476 5618 126532 5630
rect 126588 5124 126644 7308
rect 126924 6692 126980 6702
rect 126924 6598 126980 6636
rect 127148 6132 127204 20636
rect 128492 20244 128548 20254
rect 127356 19628 127620 19638
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127356 19562 127620 19572
rect 127356 18060 127620 18070
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127356 17994 127620 18004
rect 127356 16492 127620 16502
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127356 16426 127620 16436
rect 127356 14924 127620 14934
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127356 14858 127620 14868
rect 127356 13356 127620 13366
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127356 13290 127620 13300
rect 127356 11788 127620 11798
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127356 11722 127620 11732
rect 128044 11508 128100 11518
rect 127356 10220 127620 10230
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127356 10154 127620 10164
rect 127356 8652 127620 8662
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127356 8586 127620 8596
rect 127932 7362 127988 7374
rect 127932 7310 127934 7362
rect 127986 7310 127988 7362
rect 127356 7084 127620 7094
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127356 7018 127620 7028
rect 127820 6580 127876 6590
rect 127372 6466 127428 6478
rect 127372 6414 127374 6466
rect 127426 6414 127428 6466
rect 127260 6132 127316 6142
rect 127148 6130 127316 6132
rect 127148 6078 127262 6130
rect 127314 6078 127316 6130
rect 127148 6076 127316 6078
rect 126812 5796 126868 5806
rect 126812 5702 126868 5740
rect 126364 4510 126366 4562
rect 126418 4510 126420 4562
rect 126364 4498 126420 4510
rect 126476 5068 126644 5124
rect 126700 5682 126756 5694
rect 126700 5630 126702 5682
rect 126754 5630 126756 5682
rect 126028 3612 126196 3668
rect 125804 800 125860 3612
rect 126028 3332 126084 3342
rect 126028 3238 126084 3276
rect 126140 2884 126196 3612
rect 126140 2818 126196 2828
rect 126252 1204 126308 4284
rect 126364 3556 126420 3566
rect 126476 3556 126532 5068
rect 126364 3554 126532 3556
rect 126364 3502 126366 3554
rect 126418 3502 126532 3554
rect 126364 3500 126532 3502
rect 126588 4898 126644 4910
rect 126588 4846 126590 4898
rect 126642 4846 126644 4898
rect 126364 3444 126420 3500
rect 126364 3378 126420 3388
rect 126588 2436 126644 4846
rect 126700 4564 126756 5630
rect 127036 5682 127092 5694
rect 127036 5630 127038 5682
rect 127090 5630 127092 5682
rect 126812 4564 126868 4574
rect 126700 4508 126812 4564
rect 126700 4338 126756 4350
rect 126700 4286 126702 4338
rect 126754 4286 126756 4338
rect 126700 3892 126756 4286
rect 126700 3826 126756 3836
rect 126252 1138 126308 1148
rect 126364 2380 126644 2436
rect 126364 800 126420 2380
rect 126812 1540 126868 4508
rect 127036 3556 127092 5630
rect 127148 5236 127204 6076
rect 127260 6066 127316 6076
rect 127372 5682 127428 6414
rect 127372 5630 127374 5682
rect 127426 5630 127428 5682
rect 127372 5618 127428 5630
rect 127708 5908 127764 5918
rect 127708 5572 127764 5852
rect 127356 5516 127620 5526
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127708 5506 127764 5516
rect 127820 5684 127876 6524
rect 127932 6020 127988 7310
rect 128044 6690 128100 11452
rect 128492 10164 128548 20188
rect 130396 20188 130452 22092
rect 130396 20132 130564 20188
rect 129836 12740 129892 12750
rect 129276 12068 129332 12078
rect 128492 10098 128548 10108
rect 129052 10164 129108 10174
rect 128828 8034 128884 8046
rect 128828 7982 128830 8034
rect 128882 7982 128884 8034
rect 128604 7588 128660 7598
rect 128380 7362 128436 7374
rect 128380 7310 128382 7362
rect 128434 7310 128436 7362
rect 128044 6638 128046 6690
rect 128098 6638 128100 6690
rect 128044 6468 128100 6638
rect 128044 6402 128100 6412
rect 128156 6804 128212 6814
rect 128044 6132 128100 6142
rect 128156 6132 128212 6748
rect 128044 6130 128212 6132
rect 128044 6078 128046 6130
rect 128098 6078 128212 6130
rect 128044 6076 128212 6078
rect 128044 6066 128100 6076
rect 127932 5954 127988 5964
rect 128268 5908 128324 5918
rect 128268 5814 128324 5852
rect 127932 5684 127988 5694
rect 127820 5682 127988 5684
rect 127820 5630 127934 5682
rect 127986 5630 127988 5682
rect 127820 5628 127988 5630
rect 127356 5450 127620 5460
rect 127820 5348 127876 5628
rect 127932 5618 127988 5628
rect 128380 5348 128436 7310
rect 128604 6804 128660 7532
rect 128604 6690 128660 6748
rect 128604 6638 128606 6690
rect 128658 6638 128660 6690
rect 128604 6626 128660 6638
rect 127148 5170 127204 5180
rect 127596 5292 127876 5348
rect 128044 5292 128436 5348
rect 128492 6468 128548 6478
rect 127260 5124 127316 5134
rect 127260 5030 127316 5068
rect 127596 5124 127652 5292
rect 127596 5058 127652 5068
rect 127708 5122 127764 5134
rect 127932 5124 127988 5134
rect 127708 5070 127710 5122
rect 127762 5070 127764 5122
rect 127708 5012 127764 5070
rect 127708 4946 127764 4956
rect 127820 5122 127988 5124
rect 127820 5070 127934 5122
rect 127986 5070 127988 5122
rect 127820 5068 127988 5070
rect 127820 4676 127876 5068
rect 127932 5058 127988 5068
rect 127708 4620 127876 4676
rect 127036 3490 127092 3500
rect 127148 4226 127204 4238
rect 127148 4174 127150 4226
rect 127202 4174 127204 4226
rect 126812 1474 126868 1484
rect 126924 3444 126980 3454
rect 127148 3388 127204 4174
rect 127356 3948 127620 3958
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127356 3882 127620 3892
rect 127596 3780 127652 3790
rect 127260 3556 127316 3566
rect 127260 3462 127316 3500
rect 127484 3556 127540 3566
rect 126924 800 126980 3388
rect 127036 3332 127204 3388
rect 127036 3108 127092 3332
rect 127036 3042 127092 3052
rect 127484 800 127540 3500
rect 127596 3330 127652 3724
rect 127708 3388 127764 4620
rect 127932 4564 127988 4574
rect 127932 4470 127988 4508
rect 127820 4450 127876 4462
rect 127820 4398 127822 4450
rect 127874 4398 127876 4450
rect 127820 4340 127876 4398
rect 128044 4340 128100 5292
rect 128156 5124 128212 5162
rect 128156 5058 128212 5068
rect 128380 5124 128436 5134
rect 128492 5124 128548 6412
rect 128380 5122 128492 5124
rect 128380 5070 128382 5122
rect 128434 5070 128492 5122
rect 128380 5068 128492 5070
rect 128380 5058 128436 5068
rect 128492 4992 128548 5068
rect 128604 6020 128660 6030
rect 127820 4284 128044 4340
rect 128044 4274 128100 4284
rect 128156 4900 128212 4910
rect 128044 4116 128100 4126
rect 128156 4116 128212 4844
rect 128604 4228 128660 5964
rect 128044 4114 128212 4116
rect 128044 4062 128046 4114
rect 128098 4062 128212 4114
rect 128044 4060 128212 4062
rect 128492 4172 128660 4228
rect 128716 4340 128772 4350
rect 128828 4340 128884 7982
rect 128940 7362 128996 7374
rect 128940 7310 128942 7362
rect 128994 7310 128996 7362
rect 128940 6916 128996 7310
rect 128940 6850 128996 6860
rect 128940 6692 128996 6702
rect 129052 6692 129108 10108
rect 129276 7700 129332 12012
rect 128940 6690 129108 6692
rect 128940 6638 128942 6690
rect 128994 6638 129108 6690
rect 128940 6636 129108 6638
rect 129164 7644 129276 7700
rect 128940 5122 128996 6636
rect 128940 5070 128942 5122
rect 128994 5070 128996 5122
rect 128940 5058 128996 5070
rect 129052 6018 129108 6030
rect 129052 5966 129054 6018
rect 129106 5966 129108 6018
rect 129052 4452 129108 5966
rect 129164 4452 129220 7644
rect 129276 7634 129332 7644
rect 129500 7362 129556 7374
rect 129500 7310 129502 7362
rect 129554 7310 129556 7362
rect 129276 5908 129332 5918
rect 129276 5010 129332 5852
rect 129276 4958 129278 5010
rect 129330 4958 129332 5010
rect 129276 4676 129332 4958
rect 129276 4610 129332 4620
rect 129276 4452 129332 4462
rect 129164 4450 129332 4452
rect 129164 4398 129278 4450
rect 129330 4398 129332 4450
rect 129164 4396 129332 4398
rect 129052 4358 129108 4396
rect 129276 4386 129332 4396
rect 128828 4284 128996 4340
rect 128044 4050 128100 4060
rect 128044 3892 128100 3902
rect 127708 3332 127876 3388
rect 127596 3278 127598 3330
rect 127650 3278 127652 3330
rect 127596 3266 127652 3278
rect 127820 3220 127876 3332
rect 127820 2324 127876 3164
rect 127820 2258 127876 2268
rect 128044 800 128100 3836
rect 128492 3668 128548 4172
rect 128492 3554 128548 3612
rect 128492 3502 128494 3554
rect 128546 3502 128548 3554
rect 128492 3490 128548 3502
rect 128604 4004 128660 4014
rect 128156 3332 128212 3342
rect 128156 3238 128212 3276
rect 128604 800 128660 3948
rect 128716 2994 128772 4284
rect 128940 3556 128996 4284
rect 129164 4226 129220 4238
rect 129164 4174 129166 4226
rect 129218 4174 129220 4226
rect 129164 4116 129220 4174
rect 129164 4050 129220 4060
rect 129164 3668 129220 3678
rect 129052 3556 129108 3566
rect 128940 3554 129108 3556
rect 128940 3502 129054 3554
rect 129106 3502 129108 3554
rect 128940 3500 129108 3502
rect 128940 3444 128996 3500
rect 129052 3490 129108 3500
rect 128940 3378 128996 3388
rect 128716 2942 128718 2994
rect 128770 2942 128772 2994
rect 128716 2930 128772 2942
rect 129164 800 129220 3612
rect 129388 3330 129444 3342
rect 129388 3278 129390 3330
rect 129442 3278 129444 3330
rect 129388 2994 129444 3278
rect 129500 3220 129556 7310
rect 129724 6578 129780 6590
rect 129724 6526 129726 6578
rect 129778 6526 129780 6578
rect 129612 6020 129668 6030
rect 129612 3388 129668 5964
rect 129724 5684 129780 6526
rect 129836 6466 129892 12684
rect 130172 8036 130228 8046
rect 129948 7700 130004 7710
rect 129948 7606 130004 7644
rect 130060 7476 130116 7486
rect 130060 6690 130116 7420
rect 130060 6638 130062 6690
rect 130114 6638 130116 6690
rect 130060 6626 130116 6638
rect 129836 6414 129838 6466
rect 129890 6414 129892 6466
rect 129836 6402 129892 6414
rect 130060 6468 130116 6478
rect 129948 5684 130004 5694
rect 129724 5682 130004 5684
rect 129724 5630 129950 5682
rect 130002 5630 130004 5682
rect 129724 5628 130004 5630
rect 129836 4898 129892 4910
rect 129836 4846 129838 4898
rect 129890 4846 129892 4898
rect 129724 4676 129780 4686
rect 129724 3668 129780 4620
rect 129836 3892 129892 4846
rect 129948 4900 130004 5628
rect 129948 4834 130004 4844
rect 130060 5460 130116 6412
rect 130060 4676 130116 5404
rect 129948 4620 130116 4676
rect 129948 4226 130004 4620
rect 129948 4174 129950 4226
rect 130002 4174 130004 4226
rect 129948 4162 130004 4174
rect 130060 4450 130116 4462
rect 130060 4398 130062 4450
rect 130114 4398 130116 4450
rect 129836 3826 129892 3836
rect 130060 3780 130116 4398
rect 130172 4452 130228 7980
rect 130284 7700 130340 7710
rect 130284 5908 130340 7644
rect 130396 7476 130452 7486
rect 130396 6132 130452 7420
rect 130508 6580 130564 20132
rect 131740 16772 131796 115500
rect 136892 115554 136948 116398
rect 139356 116450 139636 116452
rect 139356 116398 139582 116450
rect 139634 116398 139636 116450
rect 139356 116396 139636 116398
rect 139356 115890 139412 116396
rect 139580 116386 139636 116396
rect 139356 115838 139358 115890
rect 139410 115838 139412 115890
rect 139356 115826 139412 115838
rect 140924 115780 140980 119200
rect 144060 117236 144116 119200
rect 144060 117170 144116 117180
rect 144956 117236 145012 117246
rect 144956 116562 145012 117180
rect 144956 116510 144958 116562
rect 145010 116510 145012 116562
rect 144956 116498 145012 116510
rect 145628 116564 145684 119200
rect 148764 116676 148820 119200
rect 148764 116610 148820 116620
rect 149548 116676 149604 116686
rect 145628 116498 145684 116508
rect 147532 116564 147588 116574
rect 147532 116470 147588 116508
rect 149548 116562 149604 116620
rect 149548 116510 149550 116562
rect 149602 116510 149604 116562
rect 149548 116498 149604 116510
rect 150332 116564 150388 119200
rect 153468 117012 153524 119200
rect 153468 116946 153524 116956
rect 150332 116498 150388 116508
rect 151452 116564 151508 116574
rect 151452 116470 151508 116508
rect 144284 116452 144340 116462
rect 144060 116450 144340 116452
rect 144060 116398 144286 116450
rect 144338 116398 144340 116450
rect 144060 116396 144340 116398
rect 142716 116060 142980 116070
rect 142772 116004 142820 116060
rect 142876 116004 142924 116060
rect 142716 115994 142980 116004
rect 144060 115890 144116 116396
rect 144284 116386 144340 116396
rect 146076 116452 146132 116462
rect 146076 116358 146132 116396
rect 146860 116452 146916 116462
rect 146860 116358 146916 116396
rect 148764 116450 148820 116462
rect 150780 116452 150836 116462
rect 148764 116398 148766 116450
rect 148818 116398 148820 116450
rect 144060 115838 144062 115890
rect 144114 115838 144116 115890
rect 144060 115826 144116 115838
rect 148764 115890 148820 116398
rect 148764 115838 148766 115890
rect 148818 115838 148820 115890
rect 148764 115826 148820 115838
rect 150444 116450 150836 116452
rect 150444 116398 150782 116450
rect 150834 116398 150836 116450
rect 150444 116396 150836 116398
rect 150444 115890 150500 116396
rect 150780 116386 150836 116396
rect 153468 116452 153524 116462
rect 150444 115838 150446 115890
rect 150498 115838 150500 115890
rect 140924 115714 140980 115724
rect 142044 115780 142100 115790
rect 142044 115686 142100 115724
rect 138460 115668 138516 115678
rect 138460 115574 138516 115612
rect 139132 115668 139188 115678
rect 139132 115574 139188 115612
rect 141148 115666 141204 115678
rect 141148 115614 141150 115666
rect 141202 115614 141204 115666
rect 136892 115502 136894 115554
rect 136946 115502 136948 115554
rect 133980 23940 134036 23950
rect 131740 16706 131796 16716
rect 133532 22372 133588 22382
rect 131516 15540 131572 15550
rect 130732 10612 130788 10622
rect 130620 8036 130676 8046
rect 130620 7942 130676 7980
rect 130620 6692 130676 6702
rect 130620 6598 130676 6636
rect 130508 6514 130564 6524
rect 130732 6466 130788 10556
rect 131516 8260 131572 15484
rect 131180 8204 131572 8260
rect 131068 8036 131124 8046
rect 130844 7700 130900 7710
rect 130844 7606 130900 7644
rect 130956 6916 131012 6926
rect 130732 6414 130734 6466
rect 130786 6414 130788 6466
rect 130732 6402 130788 6414
rect 130844 6692 130900 6702
rect 130396 6076 130788 6132
rect 130284 5906 130564 5908
rect 130284 5854 130286 5906
rect 130338 5854 130564 5906
rect 130284 5852 130564 5854
rect 130284 5842 130340 5852
rect 130284 5684 130340 5694
rect 130284 5682 130452 5684
rect 130284 5630 130286 5682
rect 130338 5630 130452 5682
rect 130284 5628 130452 5630
rect 130284 5618 130340 5628
rect 130284 4452 130340 4462
rect 130172 4450 130340 4452
rect 130172 4398 130286 4450
rect 130338 4398 130340 4450
rect 130172 4396 130340 4398
rect 130284 4386 130340 4396
rect 130060 3714 130116 3724
rect 130284 3892 130340 3902
rect 129948 3668 130004 3678
rect 129724 3666 130004 3668
rect 129724 3614 129950 3666
rect 130002 3614 130004 3666
rect 129724 3612 130004 3614
rect 129948 3602 130004 3612
rect 130172 3444 130228 3482
rect 129612 3332 129780 3388
rect 130172 3378 130228 3388
rect 129500 3154 129556 3164
rect 129388 2942 129390 2994
rect 129442 2942 129444 2994
rect 129388 1092 129444 2942
rect 129388 1026 129444 1036
rect 129724 800 129780 3332
rect 130060 3330 130116 3342
rect 130060 3278 130062 3330
rect 130114 3278 130116 3330
rect 130060 3220 130116 3278
rect 130060 3154 130116 3164
rect 130284 800 130340 3836
rect 130396 980 130452 5628
rect 130508 5122 130564 5852
rect 130508 5070 130510 5122
rect 130562 5070 130564 5122
rect 130508 2772 130564 5070
rect 130732 5122 130788 6076
rect 130732 5070 130734 5122
rect 130786 5070 130788 5122
rect 130620 5012 130676 5022
rect 130620 4918 130676 4956
rect 130508 2706 130564 2716
rect 130732 2324 130788 5070
rect 130844 6018 130900 6636
rect 130956 6690 131012 6860
rect 130956 6638 130958 6690
rect 131010 6638 131012 6690
rect 130956 6626 131012 6638
rect 131068 6468 131124 7980
rect 130844 5966 130846 6018
rect 130898 5966 130900 6018
rect 130844 4900 130900 5966
rect 130844 4834 130900 4844
rect 130956 6412 131124 6468
rect 130844 4676 130900 4686
rect 130844 4450 130900 4620
rect 130844 4398 130846 4450
rect 130898 4398 130900 4450
rect 130844 4386 130900 4398
rect 130732 2258 130788 2268
rect 130844 3556 130900 3566
rect 130396 924 130564 980
rect 98588 690 98644 700
rect 98896 0 99008 800
rect 99456 0 99568 800
rect 100016 0 100128 800
rect 100576 0 100688 800
rect 101136 0 101248 800
rect 101696 0 101808 800
rect 102256 0 102368 800
rect 102816 0 102928 800
rect 103376 0 103488 800
rect 103936 0 104048 800
rect 104496 0 104608 800
rect 105056 0 105168 800
rect 105616 0 105728 800
rect 106176 0 106288 800
rect 106736 0 106848 800
rect 107296 0 107408 800
rect 107856 0 107968 800
rect 108416 0 108528 800
rect 108976 0 109088 800
rect 109536 0 109648 800
rect 110096 0 110208 800
rect 110656 0 110768 800
rect 111216 0 111328 800
rect 111776 0 111888 800
rect 112336 0 112448 800
rect 112896 0 113008 800
rect 113456 0 113568 800
rect 114016 0 114128 800
rect 114576 0 114688 800
rect 115136 0 115248 800
rect 115696 0 115808 800
rect 116256 0 116368 800
rect 116816 0 116928 800
rect 117376 0 117488 800
rect 117936 0 118048 800
rect 118496 0 118608 800
rect 119056 0 119168 800
rect 119616 0 119728 800
rect 120176 0 120288 800
rect 120736 0 120848 800
rect 121296 0 121408 800
rect 121856 0 121968 800
rect 122416 0 122528 800
rect 122976 0 123088 800
rect 123536 0 123648 800
rect 124096 0 124208 800
rect 124656 0 124768 800
rect 125216 0 125328 800
rect 125776 0 125888 800
rect 126336 0 126448 800
rect 126896 0 127008 800
rect 127456 0 127568 800
rect 128016 0 128128 800
rect 128576 0 128688 800
rect 129136 0 129248 800
rect 129696 0 129808 800
rect 130256 0 130368 800
rect 130508 756 130564 924
rect 130844 800 130900 3500
rect 130956 3444 131012 6412
rect 131180 6132 131236 8204
rect 131404 8036 131460 8046
rect 131180 6018 131236 6076
rect 131180 5966 131182 6018
rect 131234 5966 131236 6018
rect 131180 5954 131236 5966
rect 131292 8034 131460 8036
rect 131292 7982 131406 8034
rect 131458 7982 131460 8034
rect 131292 7980 131460 7982
rect 131180 5124 131236 5134
rect 131068 5010 131124 5022
rect 131068 4958 131070 5010
rect 131122 4958 131124 5010
rect 131068 4788 131124 4958
rect 131068 4722 131124 4732
rect 131068 4452 131124 4462
rect 131068 4358 131124 4396
rect 131180 4226 131236 5068
rect 131180 4174 131182 4226
rect 131234 4174 131236 4226
rect 131180 4162 131236 4174
rect 131292 3668 131348 7980
rect 131404 7970 131460 7980
rect 131516 7698 131572 8204
rect 131964 8036 132020 8046
rect 131964 8034 132244 8036
rect 131964 7982 131966 8034
rect 132018 7982 132244 8034
rect 131964 7980 132244 7982
rect 131964 7970 132020 7980
rect 131516 7646 131518 7698
rect 131570 7646 131572 7698
rect 131516 7634 131572 7646
rect 131964 7476 132020 7486
rect 131964 7382 132020 7420
rect 131628 6466 131684 6478
rect 131628 6414 131630 6466
rect 131682 6414 131684 6466
rect 131628 5236 131684 6414
rect 131740 6020 131796 6030
rect 131740 5926 131796 5964
rect 132076 5684 132132 5694
rect 131292 3602 131348 3612
rect 131404 5180 131684 5236
rect 131740 5236 131796 5246
rect 130956 3378 131012 3388
rect 131180 3330 131236 3342
rect 131180 3278 131182 3330
rect 131234 3278 131236 3330
rect 131180 2548 131236 3278
rect 131180 2482 131236 2492
rect 131404 800 131460 5180
rect 131740 5142 131796 5180
rect 131628 5010 131684 5022
rect 131628 4958 131630 5010
rect 131682 4958 131684 5010
rect 131628 4564 131684 4958
rect 131852 4898 131908 4910
rect 131852 4846 131854 4898
rect 131906 4846 131908 4898
rect 131684 4508 131796 4564
rect 131628 4498 131684 4508
rect 131740 4450 131796 4508
rect 131740 4398 131742 4450
rect 131794 4398 131796 4450
rect 131740 4386 131796 4398
rect 131516 3668 131572 3678
rect 131516 3554 131572 3612
rect 131516 3502 131518 3554
rect 131570 3502 131572 3554
rect 131516 3490 131572 3502
rect 131852 3332 131908 4846
rect 131852 3266 131908 3276
rect 131964 4450 132020 4462
rect 131964 4398 131966 4450
rect 132018 4398 132020 4450
rect 131964 3220 132020 4398
rect 132076 4226 132132 5628
rect 132076 4174 132078 4226
rect 132130 4174 132132 4226
rect 132076 4162 132132 4174
rect 132188 4004 132244 7980
rect 132972 8034 133028 8046
rect 132972 7982 132974 8034
rect 133026 7982 133028 8034
rect 132412 7700 132468 7710
rect 132412 7606 132468 7644
rect 132748 7362 132804 7374
rect 132748 7310 132750 7362
rect 132802 7310 132804 7362
rect 132300 6916 132356 6926
rect 132300 6690 132356 6860
rect 132300 6638 132302 6690
rect 132354 6638 132356 6690
rect 132300 6626 132356 6638
rect 132636 6356 132692 6366
rect 132636 6018 132692 6300
rect 132636 5966 132638 6018
rect 132690 5966 132692 6018
rect 132636 5954 132692 5966
rect 132748 5348 132804 7310
rect 132748 5282 132804 5292
rect 132860 7250 132916 7262
rect 132860 7198 132862 7250
rect 132914 7198 132916 7250
rect 132188 3892 132244 3948
rect 132076 3836 132244 3892
rect 132412 4340 132468 4350
rect 132076 3554 132132 3836
rect 132076 3502 132078 3554
rect 132130 3502 132132 3554
rect 132076 3490 132132 3502
rect 132188 3668 132244 3678
rect 131964 3154 132020 3164
rect 132188 2996 132244 3612
rect 132412 3330 132468 4284
rect 132636 4340 132692 4350
rect 132860 4340 132916 7198
rect 132972 6244 133028 7982
rect 132972 6178 133028 6188
rect 133084 7700 133140 7710
rect 132972 6020 133028 6030
rect 132972 5926 133028 5964
rect 133084 5346 133140 7644
rect 133532 7700 133588 22316
rect 133756 13524 133812 13534
rect 133532 7634 133588 7644
rect 133644 8034 133700 8046
rect 133644 7982 133646 8034
rect 133698 7982 133700 8034
rect 133196 7362 133252 7374
rect 133196 7310 133198 7362
rect 133250 7310 133252 7362
rect 133196 7250 133252 7310
rect 133196 7198 133198 7250
rect 133250 7198 133252 7250
rect 133196 7186 133252 7198
rect 133644 6804 133700 7982
rect 133532 6748 133700 6804
rect 133308 6466 133364 6478
rect 133308 6414 133310 6466
rect 133362 6414 133364 6466
rect 133084 5294 133086 5346
rect 133138 5294 133140 5346
rect 133084 4676 133140 5294
rect 133196 6244 133252 6254
rect 133196 5684 133252 6188
rect 133196 5346 133252 5628
rect 133196 5294 133198 5346
rect 133250 5294 133252 5346
rect 133196 5282 133252 5294
rect 133084 4610 133140 4620
rect 132972 4452 133028 4462
rect 133196 4452 133252 4462
rect 132972 4450 133252 4452
rect 132972 4398 132974 4450
rect 133026 4398 133198 4450
rect 133250 4398 133252 4450
rect 132972 4396 133252 4398
rect 132972 4386 133028 4396
rect 133196 4386 133252 4396
rect 132636 4338 132916 4340
rect 132636 4286 132638 4338
rect 132690 4286 132916 4338
rect 132636 4284 132916 4286
rect 132636 3892 132692 4284
rect 132636 3826 132692 3836
rect 133308 3668 133364 6414
rect 133420 5348 133476 5358
rect 133420 5254 133476 5292
rect 133532 4900 133588 6748
rect 133756 6244 133812 13468
rect 133868 6468 133924 6478
rect 133868 6374 133924 6412
rect 133756 6188 133924 6244
rect 133868 6130 133924 6188
rect 133868 6078 133870 6130
rect 133922 6078 133924 6130
rect 133868 6066 133924 6078
rect 133756 6018 133812 6030
rect 133756 5966 133758 6018
rect 133810 5966 133812 6018
rect 133756 5236 133812 5966
rect 133980 5908 134036 23884
rect 135548 22484 135604 22494
rect 134764 18676 134820 18686
rect 134428 7700 134484 7710
rect 134428 7606 134484 7644
rect 133868 5852 134036 5908
rect 134092 7362 134148 7374
rect 134092 7310 134094 7362
rect 134146 7310 134148 7362
rect 133868 5460 133924 5852
rect 133980 5684 134036 5694
rect 133980 5590 134036 5628
rect 133868 5394 133924 5404
rect 133756 5180 133924 5236
rect 133644 5124 133700 5134
rect 133644 5030 133700 5068
rect 133756 5010 133812 5022
rect 133756 4958 133758 5010
rect 133810 4958 133812 5010
rect 133756 4900 133812 4958
rect 133868 5012 133924 5180
rect 133868 4946 133924 4956
rect 133980 5124 134036 5134
rect 134092 5124 134148 7310
rect 134652 7140 134708 7150
rect 134316 6466 134372 6478
rect 134316 6414 134318 6466
rect 134370 6414 134372 6466
rect 134036 5068 134148 5124
rect 134204 6356 134260 6366
rect 133532 4844 133700 4900
rect 133420 4452 133476 4462
rect 133420 4450 133588 4452
rect 133420 4398 133422 4450
rect 133474 4398 133588 4450
rect 133420 4396 133588 4398
rect 133420 4386 133476 4396
rect 133532 4338 133588 4396
rect 133532 4286 133534 4338
rect 133586 4286 133588 4338
rect 133532 4274 133588 4286
rect 133084 3612 133364 3668
rect 133420 3780 133476 3790
rect 132412 3278 132414 3330
rect 132466 3278 132468 3330
rect 132412 3266 132468 3278
rect 132524 3444 132580 3454
rect 131964 2940 132244 2996
rect 131964 800 132020 2940
rect 132524 800 132580 3388
rect 132972 3330 133028 3342
rect 132972 3278 132974 3330
rect 133026 3278 133028 3330
rect 132972 2660 133028 3278
rect 132972 2594 133028 2604
rect 133084 800 133140 3612
rect 133308 3444 133364 3454
rect 133420 3444 133476 3724
rect 133644 3556 133700 4844
rect 133756 4834 133812 4844
rect 133868 4788 133924 4798
rect 133756 4676 133812 4686
rect 133756 4562 133812 4620
rect 133756 4510 133758 4562
rect 133810 4510 133812 4562
rect 133756 4498 133812 4510
rect 133868 4450 133924 4732
rect 133980 4676 134036 5068
rect 134204 5012 134260 6300
rect 134316 6020 134372 6414
rect 134652 6130 134708 7084
rect 134764 6692 134820 18620
rect 135100 8036 135156 8046
rect 134764 6626 134820 6636
rect 134876 8034 135156 8036
rect 134876 7982 135102 8034
rect 135154 7982 135156 8034
rect 134876 7980 135156 7982
rect 134876 6132 134932 7980
rect 135100 7970 135156 7980
rect 135436 8034 135492 8046
rect 135436 7982 135438 8034
rect 135490 7982 135492 8034
rect 135436 7700 135492 7982
rect 135100 7644 135492 7700
rect 135548 7812 135604 22428
rect 135100 7140 135156 7644
rect 135212 7364 135268 7374
rect 135212 7362 135380 7364
rect 135212 7310 135214 7362
rect 135266 7310 135380 7362
rect 135212 7308 135380 7310
rect 135212 7298 135268 7308
rect 135100 7084 135268 7140
rect 134652 6078 134654 6130
rect 134706 6078 134708 6130
rect 134652 6066 134708 6078
rect 134764 6076 134932 6132
rect 134988 6466 135044 6478
rect 134988 6414 134990 6466
rect 135042 6414 135044 6466
rect 134540 6020 134596 6030
rect 134316 5964 134540 6020
rect 134540 5684 134596 5964
rect 134540 5618 134596 5628
rect 134764 5572 134820 6076
rect 134876 5908 134932 5946
rect 134876 5842 134932 5852
rect 134540 5460 134596 5470
rect 134316 5012 134372 5022
rect 134204 5010 134372 5012
rect 134204 4958 134318 5010
rect 134370 4958 134372 5010
rect 134204 4956 134372 4958
rect 134316 4946 134372 4956
rect 133980 4620 134148 4676
rect 133868 4398 133870 4450
rect 133922 4398 133924 4450
rect 133868 4386 133924 4398
rect 133868 4228 133924 4238
rect 133644 3490 133700 3500
rect 133756 3780 133812 3790
rect 133308 3442 133476 3444
rect 133308 3390 133310 3442
rect 133362 3390 133476 3442
rect 133308 3388 133476 3390
rect 133308 3378 133364 3388
rect 133756 3332 133812 3724
rect 133644 3276 133812 3332
rect 133868 3330 133924 4172
rect 133868 3278 133870 3330
rect 133922 3278 133924 3330
rect 133644 800 133700 3276
rect 133868 3266 133924 3278
rect 134092 3108 134148 4620
rect 134428 4340 134484 4378
rect 134428 4274 134484 4284
rect 134540 4226 134596 5404
rect 134652 5010 134708 5022
rect 134652 4958 134654 5010
rect 134706 4958 134708 5010
rect 134652 4788 134708 4958
rect 134652 4722 134708 4732
rect 134764 4450 134820 5516
rect 134764 4398 134766 4450
rect 134818 4398 134820 4450
rect 134764 4386 134820 4398
rect 134540 4174 134542 4226
rect 134594 4174 134596 4226
rect 134540 4162 134596 4174
rect 134316 4004 134372 4014
rect 134204 3556 134260 3566
rect 134204 3462 134260 3500
rect 134316 3332 134372 3948
rect 134988 3332 135044 6414
rect 135100 5012 135156 5022
rect 135100 3442 135156 4956
rect 135212 3668 135268 7084
rect 135324 6132 135380 7308
rect 135324 5908 135380 6076
rect 135436 5908 135492 5918
rect 135324 5906 135492 5908
rect 135324 5854 135438 5906
rect 135490 5854 135492 5906
rect 135324 5852 135492 5854
rect 135436 5348 135492 5852
rect 135548 5460 135604 7756
rect 135772 19124 135828 19134
rect 135660 7362 135716 7374
rect 135660 7310 135662 7362
rect 135714 7310 135716 7362
rect 135660 6020 135716 7310
rect 135772 6914 135828 19068
rect 136780 17780 136836 17790
rect 136668 12292 136724 12302
rect 136668 8260 136724 12236
rect 136780 8596 136836 17724
rect 136892 17668 136948 115502
rect 140700 115556 140756 115566
rect 141148 115556 141204 115614
rect 143164 115668 143220 115678
rect 143164 115574 143220 115612
rect 143836 115668 143892 115678
rect 143836 115574 143892 115612
rect 147868 115668 147924 115678
rect 147868 115574 147924 115612
rect 148540 115668 148596 115678
rect 148540 115574 148596 115612
rect 140700 115554 141204 115556
rect 140700 115502 140702 115554
rect 140754 115502 141204 115554
rect 140700 115500 141204 115502
rect 140700 19348 140756 115500
rect 142716 114492 142980 114502
rect 142772 114436 142820 114492
rect 142876 114436 142924 114492
rect 142716 114426 142980 114436
rect 142716 112924 142980 112934
rect 142772 112868 142820 112924
rect 142876 112868 142924 112924
rect 142716 112858 142980 112868
rect 142716 111356 142980 111366
rect 142772 111300 142820 111356
rect 142876 111300 142924 111356
rect 142716 111290 142980 111300
rect 142716 109788 142980 109798
rect 142772 109732 142820 109788
rect 142876 109732 142924 109788
rect 142716 109722 142980 109732
rect 142716 108220 142980 108230
rect 142772 108164 142820 108220
rect 142876 108164 142924 108220
rect 142716 108154 142980 108164
rect 142716 106652 142980 106662
rect 142772 106596 142820 106652
rect 142876 106596 142924 106652
rect 142716 106586 142980 106596
rect 142716 105084 142980 105094
rect 142772 105028 142820 105084
rect 142876 105028 142924 105084
rect 142716 105018 142980 105028
rect 142716 103516 142980 103526
rect 142772 103460 142820 103516
rect 142876 103460 142924 103516
rect 142716 103450 142980 103460
rect 142716 101948 142980 101958
rect 142772 101892 142820 101948
rect 142876 101892 142924 101948
rect 142716 101882 142980 101892
rect 142716 100380 142980 100390
rect 142772 100324 142820 100380
rect 142876 100324 142924 100380
rect 142716 100314 142980 100324
rect 142716 98812 142980 98822
rect 142772 98756 142820 98812
rect 142876 98756 142924 98812
rect 142716 98746 142980 98756
rect 142716 97244 142980 97254
rect 142772 97188 142820 97244
rect 142876 97188 142924 97244
rect 142716 97178 142980 97188
rect 142716 95676 142980 95686
rect 142772 95620 142820 95676
rect 142876 95620 142924 95676
rect 142716 95610 142980 95620
rect 142716 94108 142980 94118
rect 142772 94052 142820 94108
rect 142876 94052 142924 94108
rect 142716 94042 142980 94052
rect 142716 92540 142980 92550
rect 142772 92484 142820 92540
rect 142876 92484 142924 92540
rect 142716 92474 142980 92484
rect 142716 90972 142980 90982
rect 142772 90916 142820 90972
rect 142876 90916 142924 90972
rect 142716 90906 142980 90916
rect 142716 89404 142980 89414
rect 142772 89348 142820 89404
rect 142876 89348 142924 89404
rect 142716 89338 142980 89348
rect 142716 87836 142980 87846
rect 142772 87780 142820 87836
rect 142876 87780 142924 87836
rect 142716 87770 142980 87780
rect 142716 86268 142980 86278
rect 142772 86212 142820 86268
rect 142876 86212 142924 86268
rect 142716 86202 142980 86212
rect 142716 84700 142980 84710
rect 142772 84644 142820 84700
rect 142876 84644 142924 84700
rect 142716 84634 142980 84644
rect 142716 83132 142980 83142
rect 142772 83076 142820 83132
rect 142876 83076 142924 83132
rect 142716 83066 142980 83076
rect 142716 81564 142980 81574
rect 142772 81508 142820 81564
rect 142876 81508 142924 81564
rect 142716 81498 142980 81508
rect 142716 79996 142980 80006
rect 142772 79940 142820 79996
rect 142876 79940 142924 79996
rect 142716 79930 142980 79940
rect 142716 78428 142980 78438
rect 142772 78372 142820 78428
rect 142876 78372 142924 78428
rect 142716 78362 142980 78372
rect 142716 76860 142980 76870
rect 142772 76804 142820 76860
rect 142876 76804 142924 76860
rect 142716 76794 142980 76804
rect 142716 75292 142980 75302
rect 142772 75236 142820 75292
rect 142876 75236 142924 75292
rect 142716 75226 142980 75236
rect 142716 73724 142980 73734
rect 142772 73668 142820 73724
rect 142876 73668 142924 73724
rect 142716 73658 142980 73668
rect 142716 72156 142980 72166
rect 142772 72100 142820 72156
rect 142876 72100 142924 72156
rect 142716 72090 142980 72100
rect 142716 70588 142980 70598
rect 142772 70532 142820 70588
rect 142876 70532 142924 70588
rect 142716 70522 142980 70532
rect 142716 69020 142980 69030
rect 142772 68964 142820 69020
rect 142876 68964 142924 69020
rect 142716 68954 142980 68964
rect 142716 67452 142980 67462
rect 142772 67396 142820 67452
rect 142876 67396 142924 67452
rect 142716 67386 142980 67396
rect 142716 65884 142980 65894
rect 142772 65828 142820 65884
rect 142876 65828 142924 65884
rect 142716 65818 142980 65828
rect 142716 64316 142980 64326
rect 142772 64260 142820 64316
rect 142876 64260 142924 64316
rect 142716 64250 142980 64260
rect 142716 62748 142980 62758
rect 142772 62692 142820 62748
rect 142876 62692 142924 62748
rect 142716 62682 142980 62692
rect 142716 61180 142980 61190
rect 142772 61124 142820 61180
rect 142876 61124 142924 61180
rect 142716 61114 142980 61124
rect 142716 59612 142980 59622
rect 142772 59556 142820 59612
rect 142876 59556 142924 59612
rect 142716 59546 142980 59556
rect 142716 58044 142980 58054
rect 142772 57988 142820 58044
rect 142876 57988 142924 58044
rect 142716 57978 142980 57988
rect 142716 56476 142980 56486
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142716 56410 142980 56420
rect 142716 54908 142980 54918
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142716 54842 142980 54852
rect 142716 53340 142980 53350
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142716 53274 142980 53284
rect 142716 51772 142980 51782
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142716 51706 142980 51716
rect 142716 50204 142980 50214
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142716 50138 142980 50148
rect 142716 48636 142980 48646
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142716 48570 142980 48580
rect 142716 47068 142980 47078
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142716 47002 142980 47012
rect 142716 45500 142980 45510
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142716 45434 142980 45444
rect 142716 43932 142980 43942
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142716 43866 142980 43876
rect 142716 42364 142980 42374
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142716 42298 142980 42308
rect 142716 40796 142980 40806
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142716 40730 142980 40740
rect 142716 39228 142980 39238
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142716 39162 142980 39172
rect 142716 37660 142980 37670
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142716 37594 142980 37604
rect 142716 36092 142980 36102
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142716 36026 142980 36036
rect 142716 34524 142980 34534
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142716 34458 142980 34468
rect 142716 32956 142980 32966
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142716 32890 142980 32900
rect 142716 31388 142980 31398
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142716 31322 142980 31332
rect 142716 29820 142980 29830
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142716 29754 142980 29764
rect 142716 28252 142980 28262
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142716 28186 142980 28196
rect 142716 26684 142980 26694
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142716 26618 142980 26628
rect 142716 25116 142980 25126
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142716 25050 142980 25060
rect 142716 23548 142980 23558
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142716 23482 142980 23492
rect 142716 21980 142980 21990
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142716 21914 142980 21924
rect 142716 20412 142980 20422
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142716 20346 142980 20356
rect 140700 19282 140756 19292
rect 142716 18844 142980 18854
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142716 18778 142980 18788
rect 136892 17602 136948 17612
rect 137228 17892 137284 17902
rect 136780 8530 136836 8540
rect 137116 13972 137172 13982
rect 136668 8194 136724 8204
rect 136668 8034 136724 8046
rect 136668 7982 136670 8034
rect 136722 7982 136724 8034
rect 135772 6862 135774 6914
rect 135826 6862 135828 6914
rect 135772 6468 135828 6862
rect 136108 7362 136164 7374
rect 136108 7310 136110 7362
rect 136162 7310 136164 7362
rect 135884 6692 135940 6702
rect 135884 6598 135940 6636
rect 135996 6468 136052 6478
rect 135772 6402 135828 6412
rect 135884 6466 136052 6468
rect 135884 6414 135998 6466
rect 136050 6414 136052 6466
rect 135884 6412 136052 6414
rect 135772 6020 135828 6058
rect 135660 5964 135772 6020
rect 135772 5954 135828 5964
rect 135548 5394 135604 5404
rect 135436 5282 135492 5292
rect 135884 5124 135940 6412
rect 135996 6402 136052 6412
rect 136108 6244 136164 7310
rect 136668 7140 136724 7982
rect 136892 7362 136948 7374
rect 136892 7310 136894 7362
rect 136946 7310 136948 7362
rect 136332 7084 136724 7140
rect 136780 7250 136836 7262
rect 136780 7198 136782 7250
rect 136834 7198 136836 7250
rect 135772 5068 135940 5124
rect 135996 6188 136164 6244
rect 136220 6244 136276 6254
rect 135996 5908 136052 6188
rect 136220 6132 136276 6188
rect 135996 5122 136052 5852
rect 135996 5070 135998 5122
rect 136050 5070 136052 5122
rect 135436 5012 135492 5022
rect 135324 5010 135492 5012
rect 135324 4958 135438 5010
rect 135490 4958 135492 5010
rect 135324 4956 135492 4958
rect 135324 4788 135380 4956
rect 135436 4946 135492 4956
rect 135660 5012 135716 5022
rect 135660 4918 135716 4956
rect 135324 4562 135380 4732
rect 135324 4510 135326 4562
rect 135378 4510 135380 4562
rect 135324 4498 135380 4510
rect 135660 4564 135716 4574
rect 135660 4450 135716 4508
rect 135660 4398 135662 4450
rect 135714 4398 135716 4450
rect 135660 4386 135716 4398
rect 135212 3602 135268 3612
rect 135436 3668 135492 3678
rect 135100 3390 135102 3442
rect 135154 3390 135156 3442
rect 135100 3378 135156 3390
rect 135324 3556 135380 3566
rect 134092 2548 134148 3052
rect 134092 2482 134148 2492
rect 134204 3276 134372 3332
rect 134764 3276 135044 3332
rect 134204 800 134260 3276
rect 134764 800 134820 3276
rect 135324 800 135380 3500
rect 135436 3554 135492 3612
rect 135436 3502 135438 3554
rect 135490 3502 135492 3554
rect 135436 3490 135492 3502
rect 135772 3108 135828 5068
rect 135996 5058 136052 5070
rect 136108 6130 136276 6132
rect 136108 6078 136222 6130
rect 136274 6078 136276 6130
rect 136108 6076 136276 6078
rect 136108 5124 136164 6076
rect 136220 6066 136276 6076
rect 136332 5460 136388 7084
rect 136668 6578 136724 6590
rect 136668 6526 136670 6578
rect 136722 6526 136724 6578
rect 136668 6468 136724 6526
rect 136108 5058 136164 5068
rect 136220 5404 136388 5460
rect 136444 6412 136724 6468
rect 135884 4898 135940 4910
rect 135884 4846 135886 4898
rect 135938 4846 135940 4898
rect 135884 4788 135940 4846
rect 135884 4722 135940 4732
rect 135772 3042 135828 3052
rect 135884 4564 135940 4574
rect 135884 800 135940 4508
rect 136108 4452 136164 4462
rect 135996 3330 136052 3342
rect 135996 3278 135998 3330
rect 136050 3278 136052 3330
rect 135996 2436 136052 3278
rect 135996 2370 136052 2380
rect 136108 1652 136164 4396
rect 136220 3780 136276 5404
rect 136220 3714 136276 3724
rect 136332 3892 136388 3902
rect 136332 3444 136388 3836
rect 136332 3350 136388 3388
rect 136108 1586 136164 1596
rect 136444 800 136500 6412
rect 136668 5796 136724 5806
rect 136668 5346 136724 5740
rect 136668 5294 136670 5346
rect 136722 5294 136724 5346
rect 136668 5282 136724 5294
rect 136780 5346 136836 7198
rect 136780 5294 136782 5346
rect 136834 5294 136836 5346
rect 136668 5012 136724 5022
rect 136668 2660 136724 4956
rect 136780 4676 136836 5294
rect 136892 6692 136948 7310
rect 136892 5348 136948 6636
rect 137004 6132 137060 6142
rect 137004 6038 137060 6076
rect 137004 5348 137060 5358
rect 136892 5346 137060 5348
rect 136892 5294 137006 5346
rect 137058 5294 137060 5346
rect 136892 5292 137060 5294
rect 137004 5282 137060 5292
rect 136780 4610 136836 4620
rect 137004 4452 137060 4462
rect 137116 4452 137172 13916
rect 137228 6692 137284 17836
rect 142716 17276 142980 17286
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142716 17210 142980 17220
rect 142716 15708 142980 15718
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142716 15642 142980 15652
rect 142604 15428 142660 15438
rect 141820 13860 141876 13870
rect 141372 13748 141428 13758
rect 139132 8932 139188 8942
rect 137788 8596 137844 8606
rect 137564 8034 137620 8046
rect 137564 7982 137566 8034
rect 137618 7982 137620 8034
rect 137340 7362 137396 7374
rect 137340 7310 137342 7362
rect 137394 7310 137396 7362
rect 137340 7028 137396 7310
rect 137340 6962 137396 6972
rect 137452 7364 137508 7374
rect 137340 6692 137396 6702
rect 137228 6636 137340 6692
rect 137228 6468 137284 6478
rect 137228 6374 137284 6412
rect 137340 6244 137396 6636
rect 137228 6188 137396 6244
rect 137228 5346 137284 6188
rect 137340 5906 137396 5918
rect 137340 5854 137342 5906
rect 137394 5854 137396 5906
rect 137340 5460 137396 5854
rect 137340 5394 137396 5404
rect 137228 5294 137230 5346
rect 137282 5294 137284 5346
rect 137228 5282 137284 5294
rect 137340 5012 137396 5022
rect 137340 4918 137396 4956
rect 137004 4450 137172 4452
rect 137004 4398 137006 4450
rect 137058 4398 137172 4450
rect 137004 4396 137172 4398
rect 137004 4386 137060 4396
rect 137340 4340 137396 4350
rect 137452 4340 137508 7308
rect 137564 6804 137620 7982
rect 137788 7698 137844 8540
rect 138796 8372 138852 8382
rect 138796 8370 139076 8372
rect 138796 8318 138798 8370
rect 138850 8318 139076 8370
rect 138796 8316 139076 8318
rect 138796 8306 138852 8316
rect 138908 8148 138964 8158
rect 137788 7646 137790 7698
rect 137842 7646 137844 7698
rect 137788 7250 137844 7646
rect 137788 7198 137790 7250
rect 137842 7198 137844 7250
rect 137788 7186 137844 7198
rect 138012 7812 138068 7822
rect 138012 7364 138068 7756
rect 138796 7700 138852 7710
rect 138908 7700 138964 8092
rect 138796 7698 138964 7700
rect 138796 7646 138798 7698
rect 138850 7646 138964 7698
rect 138796 7644 138964 7646
rect 138236 7364 138292 7374
rect 138012 7362 138292 7364
rect 138012 7310 138238 7362
rect 138290 7310 138292 7362
rect 138012 7308 138292 7310
rect 137564 6738 137620 6748
rect 137676 6468 137732 6478
rect 137564 6466 137732 6468
rect 137564 6414 137678 6466
rect 137730 6414 137732 6466
rect 137564 6412 137732 6414
rect 137564 5460 137620 6412
rect 137676 6402 137732 6412
rect 137564 5394 137620 5404
rect 137676 6244 137732 6254
rect 137676 5348 137732 6188
rect 137788 5796 137844 5806
rect 137788 5702 137844 5740
rect 137340 4338 137508 4340
rect 137340 4286 137342 4338
rect 137394 4286 137508 4338
rect 137340 4284 137508 4286
rect 137564 4340 137620 4350
rect 137676 4340 137732 5292
rect 137788 5236 137844 5246
rect 137788 5142 137844 5180
rect 137900 5012 137956 5022
rect 137900 4918 137956 4956
rect 137564 4338 137732 4340
rect 137564 4286 137566 4338
rect 137618 4286 137732 4338
rect 137564 4284 137732 4286
rect 138012 4340 138068 7308
rect 138236 7298 138292 7308
rect 138796 7364 138852 7644
rect 138796 7298 138852 7308
rect 138236 7140 138292 7150
rect 138236 6804 138292 7084
rect 138124 6466 138180 6478
rect 138124 6414 138126 6466
rect 138178 6414 138180 6466
rect 138124 5908 138180 6414
rect 138124 5842 138180 5852
rect 138124 4898 138180 4910
rect 138124 4846 138126 4898
rect 138178 4846 138180 4898
rect 138124 4564 138180 4846
rect 138236 4788 138292 6748
rect 138684 6692 138740 6702
rect 138684 6466 138740 6636
rect 138684 6414 138686 6466
rect 138738 6414 138740 6466
rect 138684 6132 138740 6414
rect 138684 6066 138740 6076
rect 138348 6020 138404 6030
rect 138348 6018 138516 6020
rect 138348 5966 138350 6018
rect 138402 5966 138516 6018
rect 138348 5964 138516 5966
rect 138348 5954 138404 5964
rect 138348 5012 138404 5022
rect 138348 4918 138404 4956
rect 138236 4732 138404 4788
rect 138236 4564 138292 4574
rect 138124 4562 138292 4564
rect 138124 4510 138238 4562
rect 138290 4510 138292 4562
rect 138124 4508 138292 4510
rect 138236 4498 138292 4508
rect 138124 4340 138180 4350
rect 138012 4338 138180 4340
rect 138012 4286 138126 4338
rect 138178 4286 138180 4338
rect 138012 4284 138180 4286
rect 137340 4274 137396 4284
rect 137564 4274 137620 4284
rect 138124 4274 138180 4284
rect 138348 4338 138404 4732
rect 138348 4286 138350 4338
rect 138402 4286 138404 4338
rect 138348 4274 138404 4286
rect 137116 4228 137172 4238
rect 137116 4134 137172 4172
rect 137340 4004 137396 4014
rect 137788 4004 137844 4014
rect 137116 3780 137172 3790
rect 137116 3554 137172 3724
rect 137340 3780 137396 3948
rect 137340 3714 137396 3724
rect 137564 3948 137788 4004
rect 137116 3502 137118 3554
rect 137170 3502 137172 3554
rect 137116 3490 137172 3502
rect 137004 3444 137060 3454
rect 136892 3332 136948 3342
rect 136892 3238 136948 3276
rect 136668 2594 136724 2604
rect 137004 800 137060 3388
rect 137564 800 137620 3948
rect 137788 3938 137844 3948
rect 138012 3780 138068 3790
rect 138012 3554 138068 3724
rect 138012 3502 138014 3554
rect 138066 3502 138068 3554
rect 138012 3490 138068 3502
rect 137788 3332 137844 3342
rect 137676 3330 137844 3332
rect 137676 3278 137790 3330
rect 137842 3278 137844 3330
rect 137676 3276 137844 3278
rect 137676 980 137732 3276
rect 137788 3266 137844 3276
rect 138460 980 138516 5964
rect 138908 5794 138964 5806
rect 138908 5742 138910 5794
rect 138962 5742 138964 5794
rect 138572 5010 138628 5022
rect 138572 4958 138574 5010
rect 138626 4958 138628 5010
rect 138572 4564 138628 4958
rect 138572 4498 138628 4508
rect 138796 4900 138852 4910
rect 138684 4340 138740 4350
rect 138572 4116 138628 4126
rect 138572 4022 138628 4060
rect 137676 914 137732 924
rect 138124 924 138516 980
rect 138124 800 138180 924
rect 138684 800 138740 4284
rect 138796 4338 138852 4844
rect 138796 4286 138798 4338
rect 138850 4286 138852 4338
rect 138796 4274 138852 4286
rect 138908 3892 138964 5742
rect 138908 3826 138964 3836
rect 139020 3780 139076 8316
rect 139132 7364 139188 8876
rect 140476 8820 140532 8830
rect 139692 8034 139748 8046
rect 139692 7982 139694 8034
rect 139746 7982 139748 8034
rect 139132 7362 139300 7364
rect 139132 7310 139134 7362
rect 139186 7310 139300 7362
rect 139132 7308 139300 7310
rect 139132 7298 139188 7308
rect 139132 6580 139188 6590
rect 139132 6486 139188 6524
rect 139132 6244 139188 6254
rect 139132 5346 139188 6188
rect 139132 5294 139134 5346
rect 139186 5294 139188 5346
rect 139132 5282 139188 5294
rect 139244 5124 139300 7308
rect 139132 5068 139300 5124
rect 139356 6468 139412 6478
rect 139580 6468 139636 6478
rect 139132 4900 139188 5068
rect 139356 5010 139412 6412
rect 139356 4958 139358 5010
rect 139410 4958 139412 5010
rect 139356 4946 139412 4958
rect 139468 6466 139636 6468
rect 139468 6414 139582 6466
rect 139634 6414 139636 6466
rect 139468 6412 139636 6414
rect 139132 4834 139188 4844
rect 139244 4898 139300 4910
rect 139244 4846 139246 4898
rect 139298 4846 139300 4898
rect 139020 3554 139076 3724
rect 139020 3502 139022 3554
rect 139074 3502 139076 3554
rect 139020 3490 139076 3502
rect 139132 3444 139188 3454
rect 139132 2660 139188 3388
rect 139244 2884 139300 4846
rect 139468 4228 139524 6412
rect 139580 6402 139636 6412
rect 139692 5908 139748 7982
rect 140140 8036 140196 8046
rect 140140 8034 140308 8036
rect 140140 7982 140142 8034
rect 140194 7982 140308 8034
rect 140140 7980 140308 7982
rect 140140 7970 140196 7980
rect 140028 7364 140084 7374
rect 140028 7362 140196 7364
rect 140028 7310 140030 7362
rect 140082 7310 140196 7362
rect 140028 7308 140196 7310
rect 140028 7298 140084 7308
rect 139804 6580 139860 6590
rect 139804 6132 139860 6524
rect 140140 6580 140196 7308
rect 140140 6514 140196 6524
rect 139916 6468 139972 6478
rect 139916 6466 140084 6468
rect 139916 6414 139918 6466
rect 139970 6414 140084 6466
rect 139916 6412 140084 6414
rect 139916 6402 139972 6412
rect 140028 6244 140084 6412
rect 140028 6178 140084 6188
rect 139916 6132 139972 6142
rect 139804 6130 139972 6132
rect 139804 6078 139918 6130
rect 139970 6078 139972 6130
rect 139804 6076 139972 6078
rect 139916 6066 139972 6076
rect 139692 5852 139972 5908
rect 139804 5684 139860 5694
rect 139692 5628 139804 5684
rect 139692 5346 139748 5628
rect 139804 5552 139860 5628
rect 139692 5294 139694 5346
rect 139746 5294 139748 5346
rect 139692 5282 139748 5294
rect 139804 5122 139860 5134
rect 139804 5070 139806 5122
rect 139858 5070 139860 5122
rect 139692 4676 139748 4686
rect 139692 4562 139748 4620
rect 139692 4510 139694 4562
rect 139746 4510 139748 4562
rect 139692 4498 139748 4510
rect 139468 4162 139524 4172
rect 139580 4450 139636 4462
rect 139580 4398 139582 4450
rect 139634 4398 139636 4450
rect 139356 3332 139412 3342
rect 139580 3332 139636 4398
rect 139804 4450 139860 5070
rect 139804 4398 139806 4450
rect 139858 4398 139860 4450
rect 139804 4386 139860 4398
rect 139356 3330 139636 3332
rect 139356 3278 139358 3330
rect 139410 3278 139636 3330
rect 139356 3276 139636 3278
rect 139692 4228 139748 4238
rect 139356 3266 139412 3276
rect 139244 2818 139300 2828
rect 139132 2604 139300 2660
rect 139244 800 139300 2604
rect 139692 2436 139748 4172
rect 139916 3556 139972 5852
rect 140140 5906 140196 5918
rect 140140 5854 140142 5906
rect 140194 5854 140196 5906
rect 139916 3490 139972 3500
rect 140028 4898 140084 4910
rect 140028 4846 140030 4898
rect 140082 4846 140084 4898
rect 139916 3330 139972 3342
rect 139916 3278 139918 3330
rect 139970 3278 139972 3330
rect 139916 3108 139972 3278
rect 139916 3042 139972 3052
rect 140028 2436 140084 4846
rect 140140 3220 140196 5854
rect 140252 4340 140308 7980
rect 140476 7364 140532 8764
rect 140924 8036 140980 8046
rect 140924 8034 141092 8036
rect 140924 7982 140926 8034
rect 140978 7982 141092 8034
rect 140924 7980 141092 7982
rect 140924 7970 140980 7980
rect 141036 7476 141092 7980
rect 141036 7420 141204 7476
rect 140476 7270 140532 7308
rect 140924 7364 140980 7374
rect 140924 7362 141092 7364
rect 140924 7310 140926 7362
rect 140978 7310 141092 7362
rect 140924 7308 141092 7310
rect 140924 7298 140980 7308
rect 140924 6468 140980 6478
rect 140588 6466 140980 6468
rect 140588 6414 140926 6466
rect 140978 6414 140980 6466
rect 140588 6412 140980 6414
rect 140588 5684 140644 6412
rect 140924 6356 140980 6412
rect 140924 6290 140980 6300
rect 140700 6244 140756 6254
rect 140700 6018 140756 6188
rect 140812 6132 140868 6142
rect 141036 6132 141092 7308
rect 140812 6038 140868 6076
rect 140924 6076 141092 6132
rect 140700 5966 140702 6018
rect 140754 5966 140756 6018
rect 140700 5954 140756 5966
rect 140588 5618 140644 5628
rect 140924 5796 140980 6076
rect 140924 5010 140980 5740
rect 140924 4958 140926 5010
rect 140978 4958 140980 5010
rect 140924 4946 140980 4958
rect 141036 5906 141092 5918
rect 141036 5854 141038 5906
rect 141090 5854 141092 5906
rect 140924 4676 140980 4686
rect 140252 4274 140308 4284
rect 140364 4450 140420 4462
rect 140364 4398 140366 4450
rect 140418 4398 140420 4450
rect 140252 3556 140308 3566
rect 140252 3462 140308 3500
rect 140364 3332 140420 4398
rect 140588 4340 140644 4350
rect 140588 4246 140644 4284
rect 140364 3266 140420 3276
rect 140476 3780 140532 3790
rect 140140 3154 140196 3164
rect 140476 3108 140532 3724
rect 140812 3332 140868 3342
rect 139692 2370 139748 2380
rect 139804 2380 140084 2436
rect 140364 3052 140532 3108
rect 140700 3330 140868 3332
rect 140700 3278 140814 3330
rect 140866 3278 140868 3330
rect 140700 3276 140868 3278
rect 139804 800 139860 2380
rect 140364 800 140420 3052
rect 140700 868 140756 3276
rect 140812 3266 140868 3276
rect 140700 802 140756 812
rect 140924 800 140980 4620
rect 141036 2884 141092 5854
rect 141148 4004 141204 7420
rect 141260 6804 141316 6814
rect 141260 6690 141316 6748
rect 141260 6638 141262 6690
rect 141314 6638 141316 6690
rect 141260 6626 141316 6638
rect 141260 5012 141316 5022
rect 141260 4918 141316 4956
rect 141372 4562 141428 13692
rect 141596 7362 141652 7374
rect 141596 7310 141598 7362
rect 141650 7310 141652 7362
rect 141596 6914 141652 7310
rect 141596 6862 141598 6914
rect 141650 6862 141652 6914
rect 141596 6850 141652 6862
rect 141708 6466 141764 6478
rect 141708 6414 141710 6466
rect 141762 6414 141764 6466
rect 141708 6244 141764 6414
rect 141708 6178 141764 6188
rect 141708 6020 141764 6030
rect 141372 4510 141374 4562
rect 141426 4510 141428 4562
rect 141372 4498 141428 4510
rect 141484 6018 141764 6020
rect 141484 5966 141710 6018
rect 141762 5966 141764 6018
rect 141484 5964 141764 5966
rect 141484 4340 141540 5964
rect 141708 5954 141764 5964
rect 141820 5010 141876 13804
rect 142492 12404 142548 12414
rect 141820 4958 141822 5010
rect 141874 4958 141876 5010
rect 141820 4946 141876 4958
rect 141932 7362 141988 7374
rect 141932 7310 141934 7362
rect 141986 7310 141988 7362
rect 141148 3554 141204 3948
rect 141148 3502 141150 3554
rect 141202 3502 141204 3554
rect 141148 3490 141204 3502
rect 141260 4284 141540 4340
rect 141596 4788 141652 4798
rect 141596 4338 141652 4732
rect 141708 4564 141764 4574
rect 141708 4470 141764 4508
rect 141596 4286 141598 4338
rect 141650 4286 141652 4338
rect 141260 2996 141316 4284
rect 141596 4274 141652 4286
rect 141820 4340 141876 4350
rect 141820 4246 141876 4284
rect 141372 4114 141428 4126
rect 141372 4062 141374 4114
rect 141426 4062 141428 4114
rect 141372 3444 141428 4062
rect 141932 3444 141988 7310
rect 142156 6914 142212 6926
rect 142156 6862 142158 6914
rect 142210 6862 142212 6914
rect 142044 6692 142100 6702
rect 142044 5124 142100 6636
rect 142044 4338 142100 5068
rect 142156 5010 142212 6862
rect 142268 6466 142324 6478
rect 142268 6414 142270 6466
rect 142322 6414 142324 6466
rect 142268 6356 142324 6414
rect 142268 5236 142324 6300
rect 142380 6468 142436 6478
rect 142380 6020 142436 6412
rect 142492 6130 142548 12348
rect 142604 7364 142660 15372
rect 142716 14140 142980 14150
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142716 14074 142980 14084
rect 143724 12964 143780 12974
rect 142716 12572 142980 12582
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142716 12506 142980 12516
rect 142716 11004 142980 11014
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142716 10938 142980 10948
rect 142716 9436 142980 9446
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142716 9370 142980 9380
rect 142716 7868 142980 7878
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142716 7802 142980 7812
rect 142716 7364 142772 7374
rect 142604 7362 142772 7364
rect 142604 7310 142718 7362
rect 142770 7310 142772 7362
rect 142604 7308 142772 7310
rect 142716 6692 142772 7308
rect 143052 7362 143108 7374
rect 143052 7310 143054 7362
rect 143106 7310 143108 7362
rect 143052 6914 143108 7310
rect 143052 6862 143054 6914
rect 143106 6862 143108 6914
rect 143052 6850 143108 6862
rect 143612 7362 143668 7374
rect 143612 7310 143614 7362
rect 143666 7310 143668 7362
rect 142716 6626 142772 6636
rect 142604 6468 142660 6478
rect 142604 6374 142660 6412
rect 143052 6468 143108 6478
rect 142716 6300 142980 6310
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142716 6234 142980 6244
rect 142492 6078 142494 6130
rect 142546 6078 142548 6130
rect 142492 6066 142548 6078
rect 142380 5926 142436 5964
rect 142716 5906 142772 5918
rect 142716 5854 142718 5906
rect 142770 5854 142772 5906
rect 142716 5684 142772 5854
rect 142268 5170 142324 5180
rect 142604 5628 142716 5684
rect 142156 4958 142158 5010
rect 142210 4958 142212 5010
rect 142156 4676 142212 4958
rect 142156 4610 142212 4620
rect 142604 4564 142660 5628
rect 142716 5618 142772 5628
rect 142940 5348 142996 5358
rect 143052 5348 143108 6412
rect 143500 6466 143556 6478
rect 143500 6414 143502 6466
rect 143554 6414 143556 6466
rect 143388 6020 143444 6030
rect 142940 5346 143108 5348
rect 142940 5294 142942 5346
rect 142994 5294 143108 5346
rect 142940 5292 143108 5294
rect 143164 6018 143444 6020
rect 143164 5966 143390 6018
rect 143442 5966 143444 6018
rect 143164 5964 143444 5966
rect 142940 5282 142996 5292
rect 143052 5122 143108 5134
rect 143052 5070 143054 5122
rect 143106 5070 143108 5122
rect 142716 4732 142980 4742
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142716 4666 142980 4676
rect 143052 4564 143108 5070
rect 142604 4508 142884 4564
rect 142044 4286 142046 4338
rect 142098 4286 142100 4338
rect 142044 4274 142100 4286
rect 142828 4338 142884 4508
rect 143052 4498 143108 4508
rect 142828 4286 142830 4338
rect 142882 4286 142884 4338
rect 142828 4274 142884 4286
rect 142268 4228 142324 4238
rect 142268 4134 142324 4172
rect 143052 4228 143108 4238
rect 143052 4134 143108 4172
rect 142604 3668 142660 3678
rect 142156 3556 142212 3566
rect 142044 3444 142100 3454
rect 141372 3388 141764 3444
rect 141932 3388 142044 3444
rect 141708 3330 141764 3388
rect 142044 3350 142100 3388
rect 141708 3278 141710 3330
rect 141762 3278 141764 3330
rect 141708 3266 141764 3278
rect 142156 3220 142212 3500
rect 142044 3164 142212 3220
rect 141260 2940 141540 2996
rect 141036 2818 141092 2828
rect 141484 800 141540 2940
rect 142044 800 142100 3164
rect 142604 800 142660 3612
rect 142940 3332 142996 3370
rect 142940 3266 142996 3276
rect 142716 3164 142980 3174
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142716 3098 142980 3108
rect 143164 800 143220 5964
rect 143388 5954 143444 5964
rect 143388 5796 143444 5806
rect 143276 5122 143332 5134
rect 143276 5070 143278 5122
rect 143330 5070 143332 5122
rect 143276 4676 143332 5070
rect 143388 5010 143444 5740
rect 143388 4958 143390 5010
rect 143442 4958 143444 5010
rect 143388 4946 143444 4958
rect 143276 4610 143332 4620
rect 143500 4564 143556 6414
rect 143388 4508 143556 4564
rect 143276 4340 143332 4350
rect 143388 4340 143444 4508
rect 143276 4338 143444 4340
rect 143276 4286 143278 4338
rect 143330 4286 143444 4338
rect 143276 4284 143444 4286
rect 143276 4274 143332 4284
rect 143276 3780 143332 3790
rect 143276 3554 143332 3724
rect 143276 3502 143278 3554
rect 143330 3502 143332 3554
rect 143276 3490 143332 3502
rect 143388 1092 143444 4284
rect 143500 4338 143556 4350
rect 143500 4286 143502 4338
rect 143554 4286 143556 4338
rect 143500 4228 143556 4286
rect 143500 4162 143556 4172
rect 143612 3556 143668 7310
rect 143724 5796 143780 12908
rect 145964 12180 146020 12190
rect 143948 7700 144004 7710
rect 143724 5730 143780 5740
rect 143836 6914 143892 6926
rect 143836 6862 143838 6914
rect 143890 6862 143892 6914
rect 143724 5572 143780 5582
rect 143724 4788 143780 5516
rect 143724 4228 143780 4732
rect 143724 4162 143780 4172
rect 143836 3780 143892 6862
rect 143948 6692 144004 7644
rect 144844 7364 144900 7374
rect 144732 7362 144900 7364
rect 144732 7310 144846 7362
rect 144898 7310 144900 7362
rect 144732 7308 144900 7310
rect 143948 6690 144116 6692
rect 143948 6638 143950 6690
rect 144002 6638 144116 6690
rect 143948 6636 144116 6638
rect 143948 6626 144004 6636
rect 143948 5794 144004 5806
rect 143948 5742 143950 5794
rect 144002 5742 144004 5794
rect 143948 5684 144004 5742
rect 143948 5618 144004 5628
rect 144060 5572 144116 6636
rect 144060 5506 144116 5516
rect 144508 6466 144564 6478
rect 144508 6414 144510 6466
rect 144562 6414 144564 6466
rect 144508 6020 144564 6414
rect 143948 5348 144004 5358
rect 143948 5254 144004 5292
rect 144508 5348 144564 5964
rect 144508 5282 144564 5292
rect 144060 5124 144116 5134
rect 144060 5030 144116 5068
rect 144172 4900 144228 4910
rect 143836 3714 143892 3724
rect 143948 4898 144228 4900
rect 143948 4846 144174 4898
rect 144226 4846 144228 4898
rect 143948 4844 144228 4846
rect 143612 3490 143668 3500
rect 143388 1026 143444 1036
rect 143724 3444 143780 3454
rect 143724 800 143780 3388
rect 143836 3330 143892 3342
rect 143836 3278 143838 3330
rect 143890 3278 143892 3330
rect 143836 2884 143892 3278
rect 143948 3332 144004 4844
rect 144172 4834 144228 4844
rect 144060 4564 144116 4574
rect 144060 4470 144116 4508
rect 144172 4228 144228 4238
rect 144172 4226 144452 4228
rect 144172 4174 144174 4226
rect 144226 4174 144452 4226
rect 144172 4172 144452 4174
rect 144172 4162 144228 4172
rect 144284 4004 144340 4014
rect 144172 3556 144228 3566
rect 144172 3462 144228 3500
rect 143948 3266 144004 3276
rect 143836 2818 143892 2828
rect 144284 800 144340 3948
rect 144396 3332 144452 4172
rect 144732 3668 144788 7308
rect 144844 7298 144900 7308
rect 145404 7362 145460 7374
rect 145404 7310 145406 7362
rect 145458 7310 145460 7362
rect 145180 6916 145236 6926
rect 145068 6468 145124 6478
rect 144732 3602 144788 3612
rect 144844 6466 145124 6468
rect 144844 6414 145070 6466
rect 145122 6414 145124 6466
rect 144844 6412 145124 6414
rect 144732 3332 144788 3342
rect 144396 3330 144788 3332
rect 144396 3278 144734 3330
rect 144786 3278 144788 3330
rect 144396 3276 144788 3278
rect 144732 3266 144788 3276
rect 144844 800 144900 6412
rect 145068 6402 145124 6412
rect 144956 6132 145012 6142
rect 144956 5010 145012 6076
rect 144956 4958 144958 5010
rect 145010 4958 145012 5010
rect 144956 4946 145012 4958
rect 145180 5796 145236 6860
rect 145292 6020 145348 6030
rect 145292 5926 145348 5964
rect 145180 4900 145236 5740
rect 145292 5012 145348 5022
rect 145292 4918 145348 4956
rect 145068 4844 145236 4900
rect 145068 4788 145124 4844
rect 144956 4732 145124 4788
rect 144956 4450 145012 4732
rect 144956 4398 144958 4450
rect 145010 4398 145012 4450
rect 144956 4386 145012 4398
rect 145180 4676 145236 4686
rect 145068 4340 145124 4350
rect 145068 4246 145124 4284
rect 145180 4338 145236 4620
rect 145404 4564 145460 7310
rect 145740 6468 145796 6478
rect 145740 6020 145796 6412
rect 145516 5906 145572 5918
rect 145516 5854 145518 5906
rect 145570 5854 145572 5906
rect 145516 5012 145572 5854
rect 145516 4946 145572 4956
rect 145180 4286 145182 4338
rect 145234 4286 145236 4338
rect 145180 3780 145236 4286
rect 145180 3714 145236 3724
rect 145292 4508 145460 4564
rect 144956 3668 145012 3678
rect 144956 3554 145012 3612
rect 144956 3502 144958 3554
rect 145010 3502 145012 3554
rect 144956 3490 145012 3502
rect 145292 3444 145348 4508
rect 145516 4452 145572 4462
rect 145740 4452 145796 5964
rect 145852 4898 145908 4910
rect 145852 4846 145854 4898
rect 145906 4846 145908 4898
rect 145852 4788 145908 4846
rect 145852 4722 145908 4732
rect 145964 4564 146020 12124
rect 150444 11172 150500 115838
rect 153468 115890 153524 116396
rect 154700 116452 154756 116462
rect 154700 116358 154756 116396
rect 153468 115838 153470 115890
rect 153522 115838 153524 115890
rect 153468 115826 153524 115838
rect 155036 115892 155092 119200
rect 158172 117122 158228 119200
rect 158172 117070 158174 117122
rect 158226 117070 158228 117122
rect 158172 117058 158228 117070
rect 159292 117122 159348 117134
rect 159292 117070 159294 117122
rect 159346 117070 159348 117122
rect 155372 117012 155428 117022
rect 155372 116562 155428 116956
rect 158076 116844 158340 116854
rect 158132 116788 158180 116844
rect 158236 116788 158284 116844
rect 158076 116778 158340 116788
rect 155372 116510 155374 116562
rect 155426 116510 155428 116562
rect 155372 116498 155428 116510
rect 159292 116562 159348 117070
rect 159740 117010 159796 119200
rect 159740 116958 159742 117010
rect 159794 116958 159796 117010
rect 159740 116946 159796 116958
rect 160412 117010 160468 117022
rect 160412 116958 160414 117010
rect 160466 116958 160468 117010
rect 159292 116510 159294 116562
rect 159346 116510 159348 116562
rect 159292 116498 159348 116510
rect 158620 116452 158676 116462
rect 158172 116450 158676 116452
rect 158172 116398 158622 116450
rect 158674 116398 158676 116450
rect 158172 116396 158676 116398
rect 155260 115892 155316 115902
rect 155036 115890 155316 115892
rect 155036 115838 155262 115890
rect 155314 115838 155316 115890
rect 155036 115836 155316 115838
rect 155260 115826 155316 115836
rect 158172 115890 158228 116396
rect 158620 116386 158676 116396
rect 160412 116338 160468 116958
rect 162876 116676 162932 119200
rect 162876 116610 162932 116620
rect 163772 116676 163828 116686
rect 163772 116562 163828 116620
rect 163772 116510 163774 116562
rect 163826 116510 163828 116562
rect 163772 116498 163828 116510
rect 163100 116452 163156 116462
rect 160412 116286 160414 116338
rect 160466 116286 160468 116338
rect 160412 116274 160468 116286
rect 162876 116450 163156 116452
rect 162876 116398 163102 116450
rect 163154 116398 163156 116450
rect 162876 116396 163156 116398
rect 158172 115838 158174 115890
rect 158226 115838 158228 115890
rect 158172 115826 158228 115838
rect 162876 115890 162932 116396
rect 163100 116386 163156 116396
rect 164444 116340 164500 119200
rect 167580 117124 167636 119200
rect 167580 117058 167636 117068
rect 168476 117124 168532 117134
rect 168476 116562 168532 117068
rect 168476 116510 168478 116562
rect 168530 116510 168532 116562
rect 168476 116498 168532 116510
rect 167804 116452 167860 116462
rect 167580 116450 167860 116452
rect 167580 116398 167806 116450
rect 167858 116398 167860 116450
rect 167580 116396 167860 116398
rect 164444 116274 164500 116284
rect 164892 116340 164948 116350
rect 164892 116246 164948 116284
rect 162876 115838 162878 115890
rect 162930 115838 162932 115890
rect 162876 115826 162932 115838
rect 167580 115890 167636 116396
rect 167804 116386 167860 116396
rect 169148 116340 169204 119200
rect 172284 116676 172340 119200
rect 173852 117908 173908 119200
rect 173852 117852 174356 117908
rect 172284 116610 172340 116620
rect 173068 116676 173124 116686
rect 173068 116562 173124 116620
rect 173068 116510 173070 116562
rect 173122 116510 173124 116562
rect 173068 116498 173124 116510
rect 170940 116452 170996 116462
rect 169148 116274 169204 116284
rect 170380 116340 170436 116350
rect 170380 116246 170436 116284
rect 167580 115838 167582 115890
rect 167634 115838 167636 115890
rect 167580 115826 167636 115838
rect 170940 115890 170996 116396
rect 172284 116452 172340 116462
rect 172284 116358 172340 116396
rect 174300 116338 174356 117852
rect 174300 116286 174302 116338
rect 174354 116286 174356 116338
rect 174300 116274 174356 116286
rect 176988 116340 177044 119200
rect 177212 116340 177268 116350
rect 176988 116338 177268 116340
rect 176988 116286 177214 116338
rect 177266 116286 177268 116338
rect 176988 116284 177268 116286
rect 177212 116274 177268 116284
rect 173436 116060 173700 116070
rect 173492 116004 173540 116060
rect 173596 116004 173644 116060
rect 173436 115994 173700 116004
rect 170940 115838 170942 115890
rect 170994 115838 170996 115890
rect 170940 115826 170996 115838
rect 178108 115892 178164 115902
rect 178108 115798 178164 115836
rect 178556 115892 178612 119200
rect 178556 115826 178612 115836
rect 152124 115668 152180 115678
rect 152124 115574 152180 115612
rect 153244 115668 153300 115678
rect 153244 115574 153300 115612
rect 157276 115668 157332 115678
rect 157276 115574 157332 115612
rect 157836 115668 157892 115678
rect 157836 115574 157892 115612
rect 161980 115668 162036 115678
rect 161980 115574 162036 115612
rect 162540 115668 162596 115678
rect 162540 115574 162596 115612
rect 166684 115668 166740 115678
rect 166684 115574 166740 115612
rect 167244 115668 167300 115678
rect 167244 115574 167300 115612
rect 170044 115668 170100 115678
rect 170044 115574 170100 115612
rect 170604 115668 170660 115678
rect 170604 115574 170660 115612
rect 158076 115276 158340 115286
rect 158132 115220 158180 115276
rect 158236 115220 158284 115276
rect 158076 115210 158340 115220
rect 173436 114492 173700 114502
rect 173492 114436 173540 114492
rect 173596 114436 173644 114492
rect 173436 114426 173700 114436
rect 158076 113708 158340 113718
rect 158132 113652 158180 113708
rect 158236 113652 158284 113708
rect 158076 113642 158340 113652
rect 173436 112924 173700 112934
rect 173492 112868 173540 112924
rect 173596 112868 173644 112924
rect 173436 112858 173700 112868
rect 158076 112140 158340 112150
rect 158132 112084 158180 112140
rect 158236 112084 158284 112140
rect 158076 112074 158340 112084
rect 173436 111356 173700 111366
rect 173492 111300 173540 111356
rect 173596 111300 173644 111356
rect 173436 111290 173700 111300
rect 158076 110572 158340 110582
rect 158132 110516 158180 110572
rect 158236 110516 158284 110572
rect 158076 110506 158340 110516
rect 173436 109788 173700 109798
rect 173492 109732 173540 109788
rect 173596 109732 173644 109788
rect 173436 109722 173700 109732
rect 158076 109004 158340 109014
rect 158132 108948 158180 109004
rect 158236 108948 158284 109004
rect 158076 108938 158340 108948
rect 173436 108220 173700 108230
rect 173492 108164 173540 108220
rect 173596 108164 173644 108220
rect 173436 108154 173700 108164
rect 158076 107436 158340 107446
rect 158132 107380 158180 107436
rect 158236 107380 158284 107436
rect 158076 107370 158340 107380
rect 173436 106652 173700 106662
rect 173492 106596 173540 106652
rect 173596 106596 173644 106652
rect 173436 106586 173700 106596
rect 158076 105868 158340 105878
rect 158132 105812 158180 105868
rect 158236 105812 158284 105868
rect 158076 105802 158340 105812
rect 173436 105084 173700 105094
rect 173492 105028 173540 105084
rect 173596 105028 173644 105084
rect 173436 105018 173700 105028
rect 158076 104300 158340 104310
rect 158132 104244 158180 104300
rect 158236 104244 158284 104300
rect 158076 104234 158340 104244
rect 173436 103516 173700 103526
rect 173492 103460 173540 103516
rect 173596 103460 173644 103516
rect 173436 103450 173700 103460
rect 158076 102732 158340 102742
rect 158132 102676 158180 102732
rect 158236 102676 158284 102732
rect 158076 102666 158340 102676
rect 173436 101948 173700 101958
rect 173492 101892 173540 101948
rect 173596 101892 173644 101948
rect 173436 101882 173700 101892
rect 158076 101164 158340 101174
rect 158132 101108 158180 101164
rect 158236 101108 158284 101164
rect 158076 101098 158340 101108
rect 173436 100380 173700 100390
rect 173492 100324 173540 100380
rect 173596 100324 173644 100380
rect 173436 100314 173700 100324
rect 158076 99596 158340 99606
rect 158132 99540 158180 99596
rect 158236 99540 158284 99596
rect 158076 99530 158340 99540
rect 173436 98812 173700 98822
rect 173492 98756 173540 98812
rect 173596 98756 173644 98812
rect 173436 98746 173700 98756
rect 158076 98028 158340 98038
rect 158132 97972 158180 98028
rect 158236 97972 158284 98028
rect 158076 97962 158340 97972
rect 173436 97244 173700 97254
rect 173492 97188 173540 97244
rect 173596 97188 173644 97244
rect 173436 97178 173700 97188
rect 158076 96460 158340 96470
rect 158132 96404 158180 96460
rect 158236 96404 158284 96460
rect 158076 96394 158340 96404
rect 173436 95676 173700 95686
rect 173492 95620 173540 95676
rect 173596 95620 173644 95676
rect 173436 95610 173700 95620
rect 158076 94892 158340 94902
rect 158132 94836 158180 94892
rect 158236 94836 158284 94892
rect 158076 94826 158340 94836
rect 173436 94108 173700 94118
rect 173492 94052 173540 94108
rect 173596 94052 173644 94108
rect 173436 94042 173700 94052
rect 158076 93324 158340 93334
rect 158132 93268 158180 93324
rect 158236 93268 158284 93324
rect 158076 93258 158340 93268
rect 173436 92540 173700 92550
rect 173492 92484 173540 92540
rect 173596 92484 173644 92540
rect 173436 92474 173700 92484
rect 158076 91756 158340 91766
rect 158132 91700 158180 91756
rect 158236 91700 158284 91756
rect 158076 91690 158340 91700
rect 173436 90972 173700 90982
rect 173492 90916 173540 90972
rect 173596 90916 173644 90972
rect 173436 90906 173700 90916
rect 158076 90188 158340 90198
rect 158132 90132 158180 90188
rect 158236 90132 158284 90188
rect 158076 90122 158340 90132
rect 173436 89404 173700 89414
rect 173492 89348 173540 89404
rect 173596 89348 173644 89404
rect 173436 89338 173700 89348
rect 158076 88620 158340 88630
rect 158132 88564 158180 88620
rect 158236 88564 158284 88620
rect 158076 88554 158340 88564
rect 173436 87836 173700 87846
rect 173492 87780 173540 87836
rect 173596 87780 173644 87836
rect 173436 87770 173700 87780
rect 158076 87052 158340 87062
rect 158132 86996 158180 87052
rect 158236 86996 158284 87052
rect 158076 86986 158340 86996
rect 173436 86268 173700 86278
rect 173492 86212 173540 86268
rect 173596 86212 173644 86268
rect 173436 86202 173700 86212
rect 158076 85484 158340 85494
rect 158132 85428 158180 85484
rect 158236 85428 158284 85484
rect 158076 85418 158340 85428
rect 173436 84700 173700 84710
rect 173492 84644 173540 84700
rect 173596 84644 173644 84700
rect 173436 84634 173700 84644
rect 158076 83916 158340 83926
rect 158132 83860 158180 83916
rect 158236 83860 158284 83916
rect 158076 83850 158340 83860
rect 173436 83132 173700 83142
rect 173492 83076 173540 83132
rect 173596 83076 173644 83132
rect 173436 83066 173700 83076
rect 158076 82348 158340 82358
rect 158132 82292 158180 82348
rect 158236 82292 158284 82348
rect 158076 82282 158340 82292
rect 173436 81564 173700 81574
rect 173492 81508 173540 81564
rect 173596 81508 173644 81564
rect 173436 81498 173700 81508
rect 158076 80780 158340 80790
rect 158132 80724 158180 80780
rect 158236 80724 158284 80780
rect 158076 80714 158340 80724
rect 173436 79996 173700 80006
rect 173492 79940 173540 79996
rect 173596 79940 173644 79996
rect 173436 79930 173700 79940
rect 158076 79212 158340 79222
rect 158132 79156 158180 79212
rect 158236 79156 158284 79212
rect 158076 79146 158340 79156
rect 173436 78428 173700 78438
rect 173492 78372 173540 78428
rect 173596 78372 173644 78428
rect 173436 78362 173700 78372
rect 158076 77644 158340 77654
rect 158132 77588 158180 77644
rect 158236 77588 158284 77644
rect 158076 77578 158340 77588
rect 173436 76860 173700 76870
rect 173492 76804 173540 76860
rect 173596 76804 173644 76860
rect 173436 76794 173700 76804
rect 158076 76076 158340 76086
rect 158132 76020 158180 76076
rect 158236 76020 158284 76076
rect 158076 76010 158340 76020
rect 173436 75292 173700 75302
rect 173492 75236 173540 75292
rect 173596 75236 173644 75292
rect 173436 75226 173700 75236
rect 158076 74508 158340 74518
rect 158132 74452 158180 74508
rect 158236 74452 158284 74508
rect 158076 74442 158340 74452
rect 173436 73724 173700 73734
rect 173492 73668 173540 73724
rect 173596 73668 173644 73724
rect 173436 73658 173700 73668
rect 158076 72940 158340 72950
rect 158132 72884 158180 72940
rect 158236 72884 158284 72940
rect 158076 72874 158340 72884
rect 173436 72156 173700 72166
rect 173492 72100 173540 72156
rect 173596 72100 173644 72156
rect 173436 72090 173700 72100
rect 158076 71372 158340 71382
rect 158132 71316 158180 71372
rect 158236 71316 158284 71372
rect 158076 71306 158340 71316
rect 173436 70588 173700 70598
rect 173492 70532 173540 70588
rect 173596 70532 173644 70588
rect 173436 70522 173700 70532
rect 158076 69804 158340 69814
rect 158132 69748 158180 69804
rect 158236 69748 158284 69804
rect 158076 69738 158340 69748
rect 173436 69020 173700 69030
rect 173492 68964 173540 69020
rect 173596 68964 173644 69020
rect 173436 68954 173700 68964
rect 158076 68236 158340 68246
rect 158132 68180 158180 68236
rect 158236 68180 158284 68236
rect 158076 68170 158340 68180
rect 173436 67452 173700 67462
rect 173492 67396 173540 67452
rect 173596 67396 173644 67452
rect 173436 67386 173700 67396
rect 158076 66668 158340 66678
rect 158132 66612 158180 66668
rect 158236 66612 158284 66668
rect 158076 66602 158340 66612
rect 173436 65884 173700 65894
rect 173492 65828 173540 65884
rect 173596 65828 173644 65884
rect 173436 65818 173700 65828
rect 158076 65100 158340 65110
rect 158132 65044 158180 65100
rect 158236 65044 158284 65100
rect 158076 65034 158340 65044
rect 173436 64316 173700 64326
rect 173492 64260 173540 64316
rect 173596 64260 173644 64316
rect 173436 64250 173700 64260
rect 158076 63532 158340 63542
rect 158132 63476 158180 63532
rect 158236 63476 158284 63532
rect 158076 63466 158340 63476
rect 173436 62748 173700 62758
rect 173492 62692 173540 62748
rect 173596 62692 173644 62748
rect 173436 62682 173700 62692
rect 158076 61964 158340 61974
rect 158132 61908 158180 61964
rect 158236 61908 158284 61964
rect 158076 61898 158340 61908
rect 173436 61180 173700 61190
rect 173492 61124 173540 61180
rect 173596 61124 173644 61180
rect 173436 61114 173700 61124
rect 158076 60396 158340 60406
rect 158132 60340 158180 60396
rect 158236 60340 158284 60396
rect 158076 60330 158340 60340
rect 173436 59612 173700 59622
rect 173492 59556 173540 59612
rect 173596 59556 173644 59612
rect 173436 59546 173700 59556
rect 158076 58828 158340 58838
rect 158132 58772 158180 58828
rect 158236 58772 158284 58828
rect 158076 58762 158340 58772
rect 173436 58044 173700 58054
rect 173492 57988 173540 58044
rect 173596 57988 173644 58044
rect 173436 57978 173700 57988
rect 158076 57260 158340 57270
rect 158132 57204 158180 57260
rect 158236 57204 158284 57260
rect 158076 57194 158340 57204
rect 173436 56476 173700 56486
rect 173492 56420 173540 56476
rect 173596 56420 173644 56476
rect 173436 56410 173700 56420
rect 158076 55692 158340 55702
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158076 55626 158340 55636
rect 173436 54908 173700 54918
rect 173492 54852 173540 54908
rect 173596 54852 173644 54908
rect 173436 54842 173700 54852
rect 158076 54124 158340 54134
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158076 54058 158340 54068
rect 173436 53340 173700 53350
rect 173492 53284 173540 53340
rect 173596 53284 173644 53340
rect 173436 53274 173700 53284
rect 158076 52556 158340 52566
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158076 52490 158340 52500
rect 173436 51772 173700 51782
rect 173492 51716 173540 51772
rect 173596 51716 173644 51772
rect 173436 51706 173700 51716
rect 158076 50988 158340 50998
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158076 50922 158340 50932
rect 173436 50204 173700 50214
rect 173492 50148 173540 50204
rect 173596 50148 173644 50204
rect 173436 50138 173700 50148
rect 158076 49420 158340 49430
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158076 49354 158340 49364
rect 173436 48636 173700 48646
rect 173492 48580 173540 48636
rect 173596 48580 173644 48636
rect 173436 48570 173700 48580
rect 158076 47852 158340 47862
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158076 47786 158340 47796
rect 173436 47068 173700 47078
rect 173492 47012 173540 47068
rect 173596 47012 173644 47068
rect 173436 47002 173700 47012
rect 158076 46284 158340 46294
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158076 46218 158340 46228
rect 173436 45500 173700 45510
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173436 45434 173700 45444
rect 158076 44716 158340 44726
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158076 44650 158340 44660
rect 173436 43932 173700 43942
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173436 43866 173700 43876
rect 158076 43148 158340 43158
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158076 43082 158340 43092
rect 173436 42364 173700 42374
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173436 42298 173700 42308
rect 158076 41580 158340 41590
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158076 41514 158340 41524
rect 173436 40796 173700 40806
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173436 40730 173700 40740
rect 158076 40012 158340 40022
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158076 39946 158340 39956
rect 173436 39228 173700 39238
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173436 39162 173700 39172
rect 158076 38444 158340 38454
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158076 38378 158340 38388
rect 173436 37660 173700 37670
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173436 37594 173700 37604
rect 158076 36876 158340 36886
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158076 36810 158340 36820
rect 173436 36092 173700 36102
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173436 36026 173700 36036
rect 158076 35308 158340 35318
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158076 35242 158340 35252
rect 173436 34524 173700 34534
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173436 34458 173700 34468
rect 158076 33740 158340 33750
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158076 33674 158340 33684
rect 173436 32956 173700 32966
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173436 32890 173700 32900
rect 158076 32172 158340 32182
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158076 32106 158340 32116
rect 173436 31388 173700 31398
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173436 31322 173700 31332
rect 158076 30604 158340 30614
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158076 30538 158340 30548
rect 173436 29820 173700 29830
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173436 29754 173700 29764
rect 158076 29036 158340 29046
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158076 28970 158340 28980
rect 173436 28252 173700 28262
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173436 28186 173700 28196
rect 158076 27468 158340 27478
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158076 27402 158340 27412
rect 173436 26684 173700 26694
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173436 26618 173700 26628
rect 158076 25900 158340 25910
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158076 25834 158340 25844
rect 173436 25116 173700 25126
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173436 25050 173700 25060
rect 169148 24500 169204 24510
rect 158076 24332 158340 24342
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158076 24266 158340 24276
rect 158076 22764 158340 22774
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158076 22698 158340 22708
rect 158076 21196 158340 21206
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158076 21130 158340 21140
rect 167356 20916 167412 20926
rect 158076 19628 158340 19638
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158076 19562 158340 19572
rect 163436 18564 163492 18574
rect 158076 18060 158340 18070
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158076 17994 158340 18004
rect 158076 16492 158340 16502
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158076 16426 158340 16436
rect 158076 14924 158340 14934
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158076 14858 158340 14868
rect 161308 13636 161364 13646
rect 158076 13356 158340 13366
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158076 13290 158340 13300
rect 158076 11788 158340 11798
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158076 11722 158340 11732
rect 150444 11106 150500 11116
rect 160412 10836 160468 10846
rect 156268 10500 156324 10510
rect 148876 9044 148932 9054
rect 146300 6466 146356 6478
rect 146300 6414 146302 6466
rect 146354 6414 146356 6466
rect 146076 5794 146132 5806
rect 146076 5742 146078 5794
rect 146130 5742 146132 5794
rect 146076 5684 146132 5742
rect 146076 5618 146132 5628
rect 146188 5012 146244 5022
rect 146188 4918 146244 4956
rect 146076 4564 146132 4574
rect 145964 4562 146132 4564
rect 145964 4510 146078 4562
rect 146130 4510 146132 4562
rect 145964 4508 146132 4510
rect 146076 4498 146132 4508
rect 145516 4450 145796 4452
rect 145516 4398 145518 4450
rect 145570 4398 145796 4450
rect 145516 4396 145796 4398
rect 145516 4386 145572 4396
rect 146300 4338 146356 6414
rect 146636 6468 146692 6478
rect 146636 6374 146692 6412
rect 146972 6468 147028 6478
rect 146748 6020 146804 6030
rect 146300 4286 146302 4338
rect 146354 4286 146356 4338
rect 146300 4004 146356 4286
rect 146300 3938 146356 3948
rect 146524 6018 146804 6020
rect 146524 5966 146750 6018
rect 146802 5966 146804 6018
rect 146524 5964 146804 5966
rect 145628 3780 145684 3790
rect 145292 3378 145348 3388
rect 145404 3556 145460 3566
rect 145404 800 145460 3500
rect 145628 3442 145684 3724
rect 146076 3668 146132 3678
rect 145628 3390 145630 3442
rect 145682 3390 145684 3442
rect 145628 3378 145684 3390
rect 145964 3444 146020 3454
rect 145964 3350 146020 3388
rect 146076 3220 146132 3612
rect 145964 3164 146132 3220
rect 145964 800 146020 3164
rect 146524 800 146580 5964
rect 146748 5954 146804 5964
rect 146748 5012 146804 5022
rect 146748 4918 146804 4956
rect 146972 4450 147028 6412
rect 147084 6468 147140 6478
rect 147644 6468 147700 6478
rect 148764 6468 148820 6478
rect 147084 6466 147252 6468
rect 147084 6414 147086 6466
rect 147138 6414 147252 6466
rect 147084 6412 147252 6414
rect 147084 6402 147140 6412
rect 147084 5236 147140 5246
rect 147084 5010 147140 5180
rect 147084 4958 147086 5010
rect 147138 4958 147140 5010
rect 147084 4946 147140 4958
rect 146972 4398 146974 4450
rect 147026 4398 147028 4450
rect 146972 4386 147028 4398
rect 147196 3556 147252 6412
rect 147532 6466 147700 6468
rect 147532 6414 147646 6466
rect 147698 6414 147700 6466
rect 147532 6412 147700 6414
rect 147308 5796 147364 5806
rect 147308 5348 147364 5740
rect 147308 5282 147364 5292
rect 147308 4340 147364 4378
rect 147308 4274 147364 4284
rect 147196 3462 147252 3500
rect 147308 4114 147364 4126
rect 147308 4062 147310 4114
rect 147362 4062 147364 4114
rect 147084 3444 147140 3454
rect 146860 3332 146916 3342
rect 146860 3238 146916 3276
rect 147084 800 147140 3388
rect 147308 2660 147364 4062
rect 147532 3668 147588 6412
rect 147644 6402 147700 6412
rect 148652 6466 148820 6468
rect 148652 6414 148766 6466
rect 148818 6414 148820 6466
rect 148652 6412 148820 6414
rect 147756 5796 147812 5806
rect 148204 5796 148260 5806
rect 147644 5794 148260 5796
rect 147644 5742 147758 5794
rect 147810 5742 148206 5794
rect 148258 5742 148260 5794
rect 147644 5740 148260 5742
rect 147644 5236 147700 5740
rect 147756 5730 147812 5740
rect 148204 5730 148260 5740
rect 147644 4788 147700 5180
rect 148652 5682 148708 6412
rect 148764 6402 148820 6412
rect 148652 5630 148654 5682
rect 148706 5630 148708 5682
rect 147756 5012 147812 5022
rect 147756 4918 147812 4956
rect 147868 4900 147924 4910
rect 147868 4898 148036 4900
rect 147868 4846 147870 4898
rect 147922 4846 148036 4898
rect 147868 4844 148036 4846
rect 147868 4834 147924 4844
rect 147644 4732 147812 4788
rect 147532 3602 147588 3612
rect 147644 4564 147700 4574
rect 147308 2594 147364 2604
rect 147644 800 147700 4508
rect 147756 4452 147812 4732
rect 147868 4452 147924 4462
rect 147756 4450 147924 4452
rect 147756 4398 147870 4450
rect 147922 4398 147924 4450
rect 147756 4396 147924 4398
rect 147868 4386 147924 4396
rect 147756 3330 147812 3342
rect 147756 3278 147758 3330
rect 147810 3278 147812 3330
rect 147756 1316 147812 3278
rect 147980 3332 148036 4844
rect 148652 4788 148708 5630
rect 148092 4452 148148 4462
rect 148092 4358 148148 4396
rect 148652 4340 148708 4732
rect 148764 5794 148820 5806
rect 148764 5742 148766 5794
rect 148818 5742 148820 5794
rect 148764 4564 148820 5742
rect 148876 5010 148932 8988
rect 151340 8484 151396 8494
rect 148876 4958 148878 5010
rect 148930 4958 148932 5010
rect 148876 4946 148932 4958
rect 148988 6804 149044 6814
rect 148764 4498 148820 4508
rect 148764 4340 148820 4350
rect 148540 4338 148820 4340
rect 148540 4286 148766 4338
rect 148818 4286 148820 4338
rect 148540 4284 148820 4286
rect 148204 4116 148260 4126
rect 148204 4114 148372 4116
rect 148204 4062 148206 4114
rect 148258 4062 148372 4114
rect 148204 4060 148372 4062
rect 148204 4050 148260 4060
rect 148204 3892 148260 3902
rect 148092 3668 148148 3678
rect 148092 3554 148148 3612
rect 148092 3502 148094 3554
rect 148146 3502 148148 3554
rect 148092 3490 148148 3502
rect 147980 3266 148036 3276
rect 147756 1250 147812 1260
rect 148204 800 148260 3836
rect 148316 2548 148372 4060
rect 148540 3444 148596 4284
rect 148764 4274 148820 4284
rect 148988 4226 149044 6748
rect 149548 5908 149604 5918
rect 149100 5794 149156 5806
rect 149100 5742 149102 5794
rect 149154 5742 149156 5794
rect 149100 5682 149156 5742
rect 149100 5630 149102 5682
rect 149154 5630 149156 5682
rect 149100 5618 149156 5630
rect 149100 5122 149156 5134
rect 149100 5070 149102 5122
rect 149154 5070 149156 5122
rect 149100 4564 149156 5070
rect 149100 4498 149156 4508
rect 149100 4340 149156 4378
rect 149100 4274 149156 4284
rect 148988 4174 148990 4226
rect 149042 4174 149044 4226
rect 148988 4162 149044 4174
rect 148652 4116 148708 4126
rect 148652 3668 148708 4060
rect 148876 3780 148932 3790
rect 148764 3668 148820 3678
rect 148652 3666 148820 3668
rect 148652 3614 148766 3666
rect 148818 3614 148820 3666
rect 148652 3612 148820 3614
rect 148764 3602 148820 3612
rect 148652 3444 148708 3454
rect 148540 3442 148708 3444
rect 148540 3390 148654 3442
rect 148706 3390 148708 3442
rect 148540 3388 148708 3390
rect 148652 3378 148708 3388
rect 148316 2482 148372 2492
rect 148876 1876 148932 3724
rect 149324 3668 149380 3678
rect 148988 3556 149044 3566
rect 148988 3462 149044 3500
rect 148764 1820 148932 1876
rect 148764 800 148820 1820
rect 149324 800 149380 3612
rect 149548 3330 149604 5852
rect 149660 5796 149716 5806
rect 149996 5796 150052 5806
rect 149660 5794 149828 5796
rect 149660 5742 149662 5794
rect 149714 5742 149828 5794
rect 149660 5740 149828 5742
rect 149660 5730 149716 5740
rect 149660 4452 149716 4462
rect 149660 4358 149716 4396
rect 149772 4340 149828 5740
rect 149772 4274 149828 4284
rect 149884 5794 150052 5796
rect 149884 5742 149998 5794
rect 150050 5742 150052 5794
rect 149884 5740 150052 5742
rect 149772 4004 149828 4014
rect 149772 3668 149828 3948
rect 149772 3602 149828 3612
rect 149884 3554 149940 5740
rect 149996 5730 150052 5740
rect 149996 4900 150052 4910
rect 149996 4450 150052 4844
rect 149996 4398 149998 4450
rect 150050 4398 150052 4450
rect 149996 3780 150052 4398
rect 149996 3714 150052 3724
rect 150108 4898 150164 4910
rect 150108 4846 150110 4898
rect 150162 4846 150164 4898
rect 149884 3502 149886 3554
rect 149938 3502 149940 3554
rect 149884 3444 149940 3502
rect 149884 3378 149940 3388
rect 149548 3278 149550 3330
rect 149602 3278 149604 3330
rect 149548 3266 149604 3278
rect 150108 2436 150164 4846
rect 150668 4900 150724 4910
rect 151228 4900 151284 4910
rect 150668 4806 150724 4844
rect 151116 4898 151284 4900
rect 151116 4846 151230 4898
rect 151282 4846 151284 4898
rect 151116 4844 151284 4846
rect 150556 4450 150612 4462
rect 150556 4398 150558 4450
rect 150610 4398 150612 4450
rect 150556 3892 150612 4398
rect 150556 3826 150612 3836
rect 151004 4340 151060 4350
rect 151116 4340 151172 4844
rect 151228 4834 151284 4844
rect 151228 4564 151284 4574
rect 151340 4564 151396 8428
rect 152572 6580 152628 6590
rect 152460 5122 152516 5134
rect 152460 5070 152462 5122
rect 152514 5070 152516 5122
rect 151228 4562 151396 4564
rect 151228 4510 151230 4562
rect 151282 4510 151396 4562
rect 151228 4508 151396 4510
rect 151788 4898 151844 4910
rect 151788 4846 151790 4898
rect 151842 4846 151844 4898
rect 151228 4498 151284 4508
rect 151060 4284 151172 4340
rect 151452 4340 151508 4350
rect 149884 2380 150164 2436
rect 150444 3556 150500 3566
rect 149884 800 149940 2380
rect 150444 800 150500 3500
rect 150780 3330 150836 3342
rect 150780 3278 150782 3330
rect 150834 3278 150836 3330
rect 150780 2996 150836 3278
rect 150780 2930 150836 2940
rect 151004 800 151060 4284
rect 151452 4246 151508 4284
rect 151676 4228 151732 4238
rect 151116 4004 151172 4014
rect 151116 3780 151172 3948
rect 151116 3554 151172 3724
rect 151116 3502 151118 3554
rect 151170 3502 151172 3554
rect 151116 3490 151172 3502
rect 151676 3330 151732 4172
rect 151676 3278 151678 3330
rect 151730 3278 151732 3330
rect 151676 3266 151732 3278
rect 151788 2436 151844 4846
rect 152012 4226 152068 4238
rect 152012 4174 152014 4226
rect 152066 4174 152068 4226
rect 152012 3780 152068 4174
rect 152012 3714 152068 3724
rect 151900 3556 151956 3566
rect 151900 3462 151956 3500
rect 151564 2380 151844 2436
rect 152124 3444 152180 3454
rect 151564 800 151620 2380
rect 152124 800 152180 3388
rect 152460 3444 152516 5070
rect 152460 3378 152516 3388
rect 152572 3330 152628 6524
rect 155372 4898 155428 4910
rect 155372 4846 155374 4898
rect 155426 4846 155428 4898
rect 153468 4452 153524 4462
rect 155148 4452 155204 4462
rect 153244 4450 153524 4452
rect 153244 4398 153470 4450
rect 153522 4398 153524 4450
rect 153244 4396 153524 4398
rect 152796 4226 152852 4238
rect 152796 4174 152798 4226
rect 152850 4174 152852 4226
rect 152796 3668 152852 4174
rect 152796 3602 152852 3612
rect 152572 3278 152574 3330
rect 152626 3278 152628 3330
rect 152572 3266 152628 3278
rect 152684 3556 152740 3566
rect 152684 800 152740 3500
rect 152908 3444 152964 3454
rect 152908 3350 152964 3388
rect 153244 800 153300 4396
rect 153468 4386 153524 4396
rect 154924 4450 155204 4452
rect 154924 4398 155150 4450
rect 155202 4398 155204 4450
rect 154924 4396 155204 4398
rect 154028 4226 154084 4238
rect 154028 4174 154030 4226
rect 154082 4174 154084 4226
rect 153692 3556 153748 3566
rect 153692 3462 153748 3500
rect 154028 3556 154084 4174
rect 154588 4226 154644 4238
rect 154588 4174 154590 4226
rect 154642 4174 154644 4226
rect 154028 3490 154084 3500
rect 154364 3668 154420 3678
rect 153916 3444 153972 3454
rect 153468 3330 153524 3342
rect 153468 3278 153470 3330
rect 153522 3278 153524 3330
rect 153468 1204 153524 3278
rect 153916 2884 153972 3388
rect 153468 1138 153524 1148
rect 153804 2828 153972 2884
rect 153804 800 153860 2828
rect 154364 800 154420 3612
rect 154588 3444 154644 4174
rect 154588 3378 154644 3388
rect 154700 3332 154756 3342
rect 154700 3238 154756 3276
rect 154924 800 154980 4396
rect 155148 4386 155204 4396
rect 155372 3668 155428 4846
rect 156268 4562 156324 10444
rect 158076 10220 158340 10230
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158076 10154 158340 10164
rect 158076 8652 158340 8662
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158076 8586 158340 8596
rect 159068 8148 159124 8158
rect 158076 7084 158340 7094
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158076 7018 158340 7028
rect 158076 5516 158340 5526
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158076 5450 158340 5460
rect 156268 4510 156270 4562
rect 156322 4510 156324 4562
rect 156268 4498 156324 4510
rect 156716 4898 156772 4910
rect 156716 4846 156718 4898
rect 156770 4846 156772 4898
rect 156492 4338 156548 4350
rect 156492 4286 156494 4338
rect 156546 4286 156548 4338
rect 155820 4228 155876 4238
rect 156492 4228 156548 4286
rect 155820 4226 156548 4228
rect 155820 4174 155822 4226
rect 155874 4174 156548 4226
rect 155820 4172 156548 4174
rect 155820 4162 155876 4172
rect 155372 3602 155428 3612
rect 155820 3668 155876 3678
rect 155484 3556 155540 3566
rect 155036 3444 155092 3454
rect 155036 3350 155092 3388
rect 155484 800 155540 3500
rect 155820 3554 155876 3612
rect 155820 3502 155822 3554
rect 155874 3502 155876 3554
rect 155820 3490 155876 3502
rect 155596 3330 155652 3342
rect 155596 3278 155598 3330
rect 155650 3278 155652 3330
rect 155596 1540 155652 3278
rect 155596 1474 155652 1484
rect 156044 800 156100 4172
rect 156492 3892 156548 3902
rect 156492 3330 156548 3836
rect 156716 3556 156772 4846
rect 158396 4900 158452 4910
rect 158396 4898 158564 4900
rect 158396 4846 158398 4898
rect 158450 4846 158564 4898
rect 158396 4844 158564 4846
rect 158396 4834 158452 4844
rect 156716 3462 156772 3500
rect 157164 4450 157220 4462
rect 157164 4398 157166 4450
rect 157218 4398 157220 4450
rect 156492 3278 156494 3330
rect 156546 3278 156548 3330
rect 156492 3266 156548 3278
rect 156604 3444 156660 3454
rect 156604 800 156660 3388
rect 157164 3444 157220 4398
rect 157164 3378 157220 3388
rect 157388 4452 157444 4462
rect 157388 3442 157444 4396
rect 158396 4450 158452 4462
rect 158396 4398 158398 4450
rect 158450 4398 158452 4450
rect 157724 4228 157780 4238
rect 157388 3390 157390 3442
rect 157442 3390 157444 3442
rect 157388 3378 157444 3390
rect 157612 4226 157780 4228
rect 157612 4174 157726 4226
rect 157778 4174 157780 4226
rect 157612 4172 157780 4174
rect 157612 3554 157668 4172
rect 157724 4162 157780 4172
rect 158076 3948 158340 3958
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158076 3882 158340 3892
rect 157612 3502 157614 3554
rect 157666 3502 157668 3554
rect 157612 2548 157668 3502
rect 157164 2492 157668 2548
rect 157724 3556 157780 3566
rect 157164 800 157220 2492
rect 157724 800 157780 3500
rect 158396 2100 158452 4398
rect 158508 3556 158564 4844
rect 159068 4562 159124 8092
rect 159516 5684 159572 5694
rect 159068 4510 159070 4562
rect 159122 4510 159124 4562
rect 159068 4498 159124 4510
rect 159292 5122 159348 5134
rect 159292 5070 159294 5122
rect 159346 5070 159348 5122
rect 159180 4226 159236 4238
rect 159180 4174 159182 4226
rect 159234 4174 159236 4226
rect 158508 3490 158564 3500
rect 158956 3556 159012 3566
rect 158956 3462 159012 3500
rect 158844 3444 158900 3454
rect 158284 2044 158452 2100
rect 158620 3330 158676 3342
rect 158620 3278 158622 3330
rect 158674 3278 158676 3330
rect 158284 800 158340 2044
rect 158620 1428 158676 3278
rect 158620 1362 158676 1372
rect 158844 800 158900 3388
rect 159180 3332 159236 4174
rect 159292 3444 159348 5070
rect 159292 3378 159348 3388
rect 159404 3556 159460 3566
rect 159180 3266 159236 3276
rect 159404 800 159460 3500
rect 159516 3330 159572 5628
rect 159964 4450 160020 4462
rect 159964 4398 159966 4450
rect 160018 4398 160020 4450
rect 159852 3444 159908 3454
rect 159852 3350 159908 3388
rect 159516 3278 159518 3330
rect 159570 3278 159572 3330
rect 159516 3266 159572 3278
rect 159964 800 160020 4398
rect 160412 3330 160468 10780
rect 161084 5122 161140 5134
rect 161084 5070 161086 5122
rect 161138 5070 161140 5122
rect 161084 4340 161140 5070
rect 161308 4562 161364 13580
rect 161308 4510 161310 4562
rect 161362 4510 161364 4562
rect 161308 4498 161364 4510
rect 161420 12068 161476 12078
rect 160748 4228 160804 4238
rect 160636 4226 160804 4228
rect 160636 4174 160750 4226
rect 160802 4174 160804 4226
rect 160636 4172 160804 4174
rect 160636 3556 160692 4172
rect 160748 4162 160804 4172
rect 160636 3462 160692 3500
rect 160412 3278 160414 3330
rect 160466 3278 160468 3330
rect 160412 3266 160468 3278
rect 160524 3444 160580 3454
rect 160524 800 160580 3388
rect 161084 800 161140 4284
rect 161308 3332 161364 3342
rect 161420 3332 161476 12012
rect 161532 4900 161588 4910
rect 161532 4898 161700 4900
rect 161532 4846 161534 4898
rect 161586 4846 161700 4898
rect 161532 4844 161700 4846
rect 161532 4834 161588 4844
rect 161532 4340 161588 4350
rect 161532 4246 161588 4284
rect 161644 3554 161700 4844
rect 162204 4452 162260 4462
rect 161644 3502 161646 3554
rect 161698 3502 161700 3554
rect 161644 3444 161700 3502
rect 161644 3378 161700 3388
rect 161756 4450 162260 4452
rect 161756 4398 162206 4450
rect 162258 4398 162260 4450
rect 161756 4396 162260 4398
rect 161308 3330 161476 3332
rect 161308 3278 161310 3330
rect 161362 3278 161476 3330
rect 161308 3276 161476 3278
rect 161308 3266 161364 3276
rect 161756 2212 161812 4396
rect 162204 4386 162260 4396
rect 162764 4228 162820 4238
rect 162764 4226 162932 4228
rect 162764 4174 162766 4226
rect 162818 4174 162932 4226
rect 162764 4172 162932 4174
rect 162764 4162 162820 4172
rect 162764 3556 162820 3566
rect 161644 2156 161812 2212
rect 162204 3444 162260 3454
rect 161644 800 161700 2156
rect 162204 800 162260 3388
rect 162540 3330 162596 3342
rect 162540 3278 162542 3330
rect 162594 3278 162596 3330
rect 162540 2324 162596 3278
rect 162540 2258 162596 2268
rect 162764 800 162820 3500
rect 162876 3444 162932 4172
rect 162876 3350 162932 3388
rect 163436 3330 163492 18508
rect 164332 7588 164388 7598
rect 163436 3278 163438 3330
rect 163490 3278 163492 3330
rect 163436 3266 163492 3278
rect 163548 4450 163604 4462
rect 163548 4398 163550 4450
rect 163602 4398 163604 4450
rect 163548 1428 163604 4398
rect 164108 4226 164164 4238
rect 164108 4174 164110 4226
rect 164162 4174 164164 4226
rect 163660 3556 163716 3566
rect 163660 3462 163716 3500
rect 164108 3556 164164 4174
rect 164108 3490 164164 3500
rect 163324 1372 163604 1428
rect 163884 3444 163940 3454
rect 163324 800 163380 1372
rect 163884 800 163940 3388
rect 164332 3330 164388 7532
rect 167132 4898 167188 4910
rect 167132 4846 167134 4898
rect 167186 4846 167188 4898
rect 165228 4452 165284 4462
rect 166908 4452 166964 4462
rect 165004 4450 165284 4452
rect 165004 4398 165230 4450
rect 165282 4398 165284 4450
rect 165004 4396 165284 4398
rect 164556 4228 164612 4238
rect 164556 4226 164724 4228
rect 164556 4174 164558 4226
rect 164610 4174 164724 4226
rect 164556 4172 164724 4174
rect 164556 4162 164612 4172
rect 164332 3278 164334 3330
rect 164386 3278 164388 3330
rect 164332 3266 164388 3278
rect 164444 3556 164500 3566
rect 164444 800 164500 3500
rect 164668 3444 164724 4172
rect 164668 3350 164724 3388
rect 165004 800 165060 4396
rect 165228 4386 165284 4396
rect 166684 4450 166964 4452
rect 166684 4398 166910 4450
rect 166962 4398 166964 4450
rect 166684 4396 166964 4398
rect 165788 4226 165844 4238
rect 165788 4174 165790 4226
rect 165842 4174 165844 4226
rect 165452 3556 165508 3566
rect 165452 3462 165508 3500
rect 165788 3556 165844 4174
rect 166348 4226 166404 4238
rect 166348 4174 166350 4226
rect 166402 4174 166404 4226
rect 165788 3490 165844 3500
rect 166124 3556 166180 3566
rect 165676 3444 165732 3454
rect 165228 3332 165284 3342
rect 165228 3238 165284 3276
rect 165676 2884 165732 3388
rect 165564 2828 165732 2884
rect 165564 800 165620 2828
rect 166124 800 166180 3500
rect 166348 3444 166404 4174
rect 166348 3378 166404 3388
rect 166460 3330 166516 3342
rect 166460 3278 166462 3330
rect 166514 3278 166516 3330
rect 166460 2436 166516 3278
rect 166460 2370 166516 2380
rect 166684 800 166740 4396
rect 166908 4386 166964 4396
rect 167132 3556 167188 4846
rect 167132 3490 167188 3500
rect 166796 3444 166852 3454
rect 166796 3350 166852 3388
rect 167244 3444 167300 3454
rect 167244 800 167300 3388
rect 167356 3330 167412 20860
rect 169148 20188 169204 24444
rect 173436 23548 173700 23558
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173436 23482 173700 23492
rect 173436 21980 173700 21990
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173436 21914 173700 21924
rect 173436 20412 173700 20422
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173436 20346 173700 20356
rect 169148 20132 169316 20188
rect 168028 4900 168084 4910
rect 168028 4898 168196 4900
rect 168028 4846 168030 4898
rect 168082 4846 168196 4898
rect 168028 4844 168196 4846
rect 168028 4834 168084 4844
rect 168028 4450 168084 4462
rect 168028 4398 168030 4450
rect 168082 4398 168084 4450
rect 167804 3668 167860 3678
rect 167580 3556 167636 3566
rect 167580 3462 167636 3500
rect 167356 3278 167358 3330
rect 167410 3278 167412 3330
rect 167356 3266 167412 3278
rect 167804 800 167860 3612
rect 168028 2324 168084 4398
rect 168140 3444 168196 4844
rect 168924 4898 168980 4910
rect 168924 4846 168926 4898
rect 168978 4846 168980 4898
rect 168924 4676 168980 4846
rect 169260 4900 169316 20132
rect 173436 18844 173700 18854
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173436 18778 173700 18788
rect 173436 17276 173700 17286
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173436 17210 173700 17220
rect 173436 15708 173700 15718
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173436 15642 173700 15652
rect 173436 14140 173700 14150
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173436 14074 173700 14084
rect 173436 12572 173700 12582
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173436 12506 173700 12516
rect 170380 11956 170436 11966
rect 169260 4834 169316 4844
rect 169372 4900 169428 4910
rect 169372 4898 169540 4900
rect 169372 4846 169374 4898
rect 169426 4846 169540 4898
rect 169372 4844 169540 4846
rect 169372 4834 169428 4844
rect 168924 4620 169428 4676
rect 169148 4452 169204 4462
rect 169036 4450 169204 4452
rect 169036 4398 169150 4450
rect 169202 4398 169204 4450
rect 169036 4396 169204 4398
rect 168140 3378 168196 3388
rect 168588 3444 168644 3454
rect 168588 3350 168644 3388
rect 168252 3330 168308 3342
rect 168252 3278 168254 3330
rect 168306 3278 168308 3330
rect 168252 2772 168308 3278
rect 168252 2706 168308 2716
rect 168028 2268 168420 2324
rect 168364 800 168420 2268
rect 169036 1652 169092 4396
rect 169148 4386 169204 4396
rect 169260 4452 169316 4462
rect 169148 3332 169204 3342
rect 169260 3332 169316 4396
rect 169148 3330 169316 3332
rect 169148 3278 169150 3330
rect 169202 3278 169316 3330
rect 169148 3276 169316 3278
rect 169372 4338 169428 4620
rect 169372 4286 169374 4338
rect 169426 4286 169428 4338
rect 169148 3266 169204 3276
rect 169036 1586 169092 1596
rect 169372 1428 169428 4286
rect 169484 3668 169540 4844
rect 170268 4452 170324 4462
rect 169484 3554 169540 3612
rect 170044 4450 170324 4452
rect 170044 4398 170270 4450
rect 170322 4398 170324 4450
rect 170044 4396 170324 4398
rect 169484 3502 169486 3554
rect 169538 3502 169540 3554
rect 169484 3490 169540 3502
rect 169596 3556 169652 3566
rect 169596 2884 169652 3500
rect 168924 1372 169428 1428
rect 169484 2828 169652 2884
rect 168924 800 168980 1372
rect 169484 800 169540 2828
rect 170044 800 170100 4396
rect 170268 4386 170324 4396
rect 170380 3330 170436 11900
rect 173436 11004 173700 11014
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173436 10938 173700 10948
rect 172172 10388 172228 10398
rect 171276 8036 171332 8046
rect 170828 4228 170884 4238
rect 170716 4226 170884 4228
rect 170716 4174 170830 4226
rect 170882 4174 170884 4226
rect 170716 4172 170884 4174
rect 170716 3556 170772 4172
rect 170828 4162 170884 4172
rect 170716 3462 170772 3500
rect 171164 3556 171220 3566
rect 170380 3278 170382 3330
rect 170434 3278 170436 3330
rect 170380 3266 170436 3278
rect 170604 3444 170660 3454
rect 170604 800 170660 3388
rect 171164 800 171220 3500
rect 171276 3330 171332 7980
rect 171948 4452 172004 4462
rect 171724 4450 172004 4452
rect 171724 4398 171950 4450
rect 172002 4398 172004 4450
rect 171724 4396 172004 4398
rect 171388 4226 171444 4238
rect 171388 4174 171390 4226
rect 171442 4174 171444 4226
rect 171388 3444 171444 4174
rect 171388 3378 171444 3388
rect 171612 3444 171668 3454
rect 171612 3350 171668 3388
rect 171276 3278 171278 3330
rect 171330 3278 171332 3330
rect 171276 3266 171332 3278
rect 171724 800 171780 4396
rect 171948 4386 172004 4396
rect 172172 3330 172228 10332
rect 173436 9436 173700 9446
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173436 9370 173700 9380
rect 173436 7868 173700 7878
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173436 7802 173700 7812
rect 173436 6300 173700 6310
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173436 6234 173700 6244
rect 173180 5348 173236 5358
rect 173068 4452 173124 4462
rect 172844 4450 173124 4452
rect 172844 4398 173070 4450
rect 173122 4398 173124 4450
rect 172844 4396 173124 4398
rect 172508 4228 172564 4238
rect 172396 4226 172564 4228
rect 172396 4174 172510 4226
rect 172562 4174 172564 4226
rect 172396 4172 172564 4174
rect 172396 3556 172452 4172
rect 172508 4162 172564 4172
rect 172396 3462 172452 3500
rect 172172 3278 172174 3330
rect 172226 3278 172228 3330
rect 172172 3266 172228 3278
rect 172284 3444 172340 3454
rect 172284 800 172340 3388
rect 172844 800 172900 4396
rect 173068 4386 173124 4396
rect 173068 3332 173124 3342
rect 173180 3332 173236 5292
rect 173436 4732 173700 4742
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173436 4666 173700 4676
rect 173628 4228 173684 4238
rect 173404 4226 173684 4228
rect 173404 4174 173630 4226
rect 173682 4174 173684 4226
rect 173404 4172 173684 4174
rect 173404 3554 173460 4172
rect 173628 4162 173684 4172
rect 173404 3502 173406 3554
rect 173458 3502 173460 3554
rect 173404 3444 173460 3502
rect 173404 3378 173460 3388
rect 173068 3330 173236 3332
rect 173068 3278 173070 3330
rect 173122 3278 173236 3330
rect 173068 3276 173236 3278
rect 173964 3332 174020 3342
rect 173068 3266 173124 3276
rect 173436 3164 173700 3174
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173436 3098 173700 3108
rect 173404 1762 173460 1774
rect 173404 1710 173406 1762
rect 173458 1710 173460 1762
rect 173404 800 173460 1710
rect 173964 800 174020 3276
rect 174300 3330 174356 3342
rect 174300 3278 174302 3330
rect 174354 3278 174356 3330
rect 174300 1762 174356 3278
rect 174972 3332 175028 3342
rect 174972 3238 175028 3276
rect 174300 1710 174302 1762
rect 174354 1710 174356 1762
rect 174300 1698 174356 1710
rect 130508 690 130564 700
rect 130816 0 130928 800
rect 131376 0 131488 800
rect 131936 0 132048 800
rect 132496 0 132608 800
rect 133056 0 133168 800
rect 133616 0 133728 800
rect 134176 0 134288 800
rect 134736 0 134848 800
rect 135296 0 135408 800
rect 135856 0 135968 800
rect 136416 0 136528 800
rect 136976 0 137088 800
rect 137536 0 137648 800
rect 138096 0 138208 800
rect 138656 0 138768 800
rect 139216 0 139328 800
rect 139776 0 139888 800
rect 140336 0 140448 800
rect 140896 0 141008 800
rect 141456 0 141568 800
rect 142016 0 142128 800
rect 142576 0 142688 800
rect 143136 0 143248 800
rect 143696 0 143808 800
rect 144256 0 144368 800
rect 144816 0 144928 800
rect 145376 0 145488 800
rect 145936 0 146048 800
rect 146496 0 146608 800
rect 147056 0 147168 800
rect 147616 0 147728 800
rect 148176 0 148288 800
rect 148736 0 148848 800
rect 149296 0 149408 800
rect 149856 0 149968 800
rect 150416 0 150528 800
rect 150976 0 151088 800
rect 151536 0 151648 800
rect 152096 0 152208 800
rect 152656 0 152768 800
rect 153216 0 153328 800
rect 153776 0 153888 800
rect 154336 0 154448 800
rect 154896 0 155008 800
rect 155456 0 155568 800
rect 156016 0 156128 800
rect 156576 0 156688 800
rect 157136 0 157248 800
rect 157696 0 157808 800
rect 158256 0 158368 800
rect 158816 0 158928 800
rect 159376 0 159488 800
rect 159936 0 160048 800
rect 160496 0 160608 800
rect 161056 0 161168 800
rect 161616 0 161728 800
rect 162176 0 162288 800
rect 162736 0 162848 800
rect 163296 0 163408 800
rect 163856 0 163968 800
rect 164416 0 164528 800
rect 164976 0 165088 800
rect 165536 0 165648 800
rect 166096 0 166208 800
rect 166656 0 166768 800
rect 167216 0 167328 800
rect 167776 0 167888 800
rect 168336 0 168448 800
rect 168896 0 169008 800
rect 169456 0 169568 800
rect 170016 0 170128 800
rect 170576 0 170688 800
rect 171136 0 171248 800
rect 171696 0 171808 800
rect 172256 0 172368 800
rect 172816 0 172928 800
rect 173376 0 173488 800
rect 173936 0 174048 800
<< via2 >>
rect 4508 116956 4564 117012
rect 5964 116956 6020 117012
rect 4476 116842 4532 116844
rect 4476 116790 4478 116842
rect 4478 116790 4530 116842
rect 4530 116790 4532 116842
rect 4476 116788 4532 116790
rect 4580 116842 4636 116844
rect 4580 116790 4582 116842
rect 4582 116790 4634 116842
rect 4634 116790 4636 116842
rect 4580 116788 4636 116790
rect 4684 116842 4740 116844
rect 4684 116790 4686 116842
rect 4686 116790 4738 116842
rect 4738 116790 4740 116842
rect 4684 116788 4740 116790
rect 2940 116508 2996 116564
rect 3388 116562 3444 116564
rect 3388 116510 3390 116562
rect 3390 116510 3442 116562
rect 3442 116510 3444 116562
rect 3388 116508 3444 116510
rect 7644 116620 7700 116676
rect 8428 116620 8484 116676
rect 9212 116508 9268 116564
rect 10108 116562 10164 116564
rect 10108 116510 10110 116562
rect 10110 116510 10162 116562
rect 10162 116510 10164 116562
rect 10108 116508 10164 116510
rect 5180 115666 5236 115668
rect 5180 115614 5182 115666
rect 5182 115614 5234 115666
rect 5234 115614 5236 115666
rect 5180 115612 5236 115614
rect 10892 116172 10948 116228
rect 11340 116226 11396 116228
rect 11340 116174 11342 116226
rect 11342 116174 11394 116226
rect 11394 116174 11396 116226
rect 11340 116172 11396 116174
rect 12348 115836 12404 115892
rect 12684 116172 12740 116228
rect 7196 115666 7252 115668
rect 7196 115614 7198 115666
rect 7198 115614 7250 115666
rect 7250 115614 7252 115666
rect 7196 115612 7252 115614
rect 7980 115666 8036 115668
rect 7980 115614 7982 115666
rect 7982 115614 8034 115666
rect 8034 115614 8036 115666
rect 7980 115612 8036 115614
rect 4476 115274 4532 115276
rect 4476 115222 4478 115274
rect 4478 115222 4530 115274
rect 4530 115222 4532 115274
rect 4476 115220 4532 115222
rect 4580 115274 4636 115276
rect 4580 115222 4582 115274
rect 4582 115222 4634 115274
rect 4634 115222 4636 115274
rect 4580 115220 4636 115222
rect 4684 115274 4740 115276
rect 4684 115222 4686 115274
rect 4686 115222 4738 115274
rect 4738 115222 4740 115274
rect 4684 115220 4740 115222
rect 4476 113706 4532 113708
rect 4476 113654 4478 113706
rect 4478 113654 4530 113706
rect 4530 113654 4532 113706
rect 4476 113652 4532 113654
rect 4580 113706 4636 113708
rect 4580 113654 4582 113706
rect 4582 113654 4634 113706
rect 4634 113654 4636 113706
rect 4580 113652 4636 113654
rect 4684 113706 4740 113708
rect 4684 113654 4686 113706
rect 4686 113654 4738 113706
rect 4738 113654 4740 113706
rect 4684 113652 4740 113654
rect 4476 112138 4532 112140
rect 4476 112086 4478 112138
rect 4478 112086 4530 112138
rect 4530 112086 4532 112138
rect 4476 112084 4532 112086
rect 4580 112138 4636 112140
rect 4580 112086 4582 112138
rect 4582 112086 4634 112138
rect 4634 112086 4636 112138
rect 4580 112084 4636 112086
rect 4684 112138 4740 112140
rect 4684 112086 4686 112138
rect 4686 112086 4738 112138
rect 4738 112086 4740 112138
rect 4684 112084 4740 112086
rect 4476 110570 4532 110572
rect 4476 110518 4478 110570
rect 4478 110518 4530 110570
rect 4530 110518 4532 110570
rect 4476 110516 4532 110518
rect 4580 110570 4636 110572
rect 4580 110518 4582 110570
rect 4582 110518 4634 110570
rect 4634 110518 4636 110570
rect 4580 110516 4636 110518
rect 4684 110570 4740 110572
rect 4684 110518 4686 110570
rect 4686 110518 4738 110570
rect 4738 110518 4740 110570
rect 4684 110516 4740 110518
rect 4476 109002 4532 109004
rect 4476 108950 4478 109002
rect 4478 108950 4530 109002
rect 4530 108950 4532 109002
rect 4476 108948 4532 108950
rect 4580 109002 4636 109004
rect 4580 108950 4582 109002
rect 4582 108950 4634 109002
rect 4634 108950 4636 109002
rect 4580 108948 4636 108950
rect 4684 109002 4740 109004
rect 4684 108950 4686 109002
rect 4686 108950 4738 109002
rect 4738 108950 4740 109002
rect 4684 108948 4740 108950
rect 11116 115666 11172 115668
rect 11116 115614 11118 115666
rect 11118 115614 11170 115666
rect 11170 115614 11172 115666
rect 11116 115612 11172 115614
rect 11676 115666 11732 115668
rect 11676 115614 11678 115666
rect 11678 115614 11730 115666
rect 11730 115614 11732 115666
rect 11676 115612 11732 115614
rect 6636 108332 6692 108388
rect 4476 107434 4532 107436
rect 4476 107382 4478 107434
rect 4478 107382 4530 107434
rect 4530 107382 4532 107434
rect 4476 107380 4532 107382
rect 4580 107434 4636 107436
rect 4580 107382 4582 107434
rect 4582 107382 4634 107434
rect 4634 107382 4636 107434
rect 4580 107380 4636 107382
rect 4684 107434 4740 107436
rect 4684 107382 4686 107434
rect 4686 107382 4738 107434
rect 4738 107382 4740 107434
rect 4684 107380 4740 107382
rect 4476 105866 4532 105868
rect 4476 105814 4478 105866
rect 4478 105814 4530 105866
rect 4530 105814 4532 105866
rect 4476 105812 4532 105814
rect 4580 105866 4636 105868
rect 4580 105814 4582 105866
rect 4582 105814 4634 105866
rect 4634 105814 4636 105866
rect 4580 105812 4636 105814
rect 4684 105866 4740 105868
rect 4684 105814 4686 105866
rect 4686 105814 4738 105866
rect 4738 105814 4740 105866
rect 4684 105812 4740 105814
rect 4476 104298 4532 104300
rect 4476 104246 4478 104298
rect 4478 104246 4530 104298
rect 4530 104246 4532 104298
rect 4476 104244 4532 104246
rect 4580 104298 4636 104300
rect 4580 104246 4582 104298
rect 4582 104246 4634 104298
rect 4634 104246 4636 104298
rect 4580 104244 4636 104246
rect 4684 104298 4740 104300
rect 4684 104246 4686 104298
rect 4686 104246 4738 104298
rect 4738 104246 4740 104298
rect 4684 104244 4740 104246
rect 4476 102730 4532 102732
rect 4476 102678 4478 102730
rect 4478 102678 4530 102730
rect 4530 102678 4532 102730
rect 4476 102676 4532 102678
rect 4580 102730 4636 102732
rect 4580 102678 4582 102730
rect 4582 102678 4634 102730
rect 4634 102678 4636 102730
rect 4580 102676 4636 102678
rect 4684 102730 4740 102732
rect 4684 102678 4686 102730
rect 4686 102678 4738 102730
rect 4738 102678 4740 102730
rect 4684 102676 4740 102678
rect 4476 101162 4532 101164
rect 4476 101110 4478 101162
rect 4478 101110 4530 101162
rect 4530 101110 4532 101162
rect 4476 101108 4532 101110
rect 4580 101162 4636 101164
rect 4580 101110 4582 101162
rect 4582 101110 4634 101162
rect 4634 101110 4636 101162
rect 4580 101108 4636 101110
rect 4684 101162 4740 101164
rect 4684 101110 4686 101162
rect 4686 101110 4738 101162
rect 4738 101110 4740 101162
rect 4684 101108 4740 101110
rect 4476 99594 4532 99596
rect 4476 99542 4478 99594
rect 4478 99542 4530 99594
rect 4530 99542 4532 99594
rect 4476 99540 4532 99542
rect 4580 99594 4636 99596
rect 4580 99542 4582 99594
rect 4582 99542 4634 99594
rect 4634 99542 4636 99594
rect 4580 99540 4636 99542
rect 4684 99594 4740 99596
rect 4684 99542 4686 99594
rect 4686 99542 4738 99594
rect 4738 99542 4740 99594
rect 4684 99540 4740 99542
rect 4476 98026 4532 98028
rect 4476 97974 4478 98026
rect 4478 97974 4530 98026
rect 4530 97974 4532 98026
rect 4476 97972 4532 97974
rect 4580 98026 4636 98028
rect 4580 97974 4582 98026
rect 4582 97974 4634 98026
rect 4634 97974 4636 98026
rect 4580 97972 4636 97974
rect 4684 98026 4740 98028
rect 4684 97974 4686 98026
rect 4686 97974 4738 98026
rect 4738 97974 4740 98026
rect 4684 97972 4740 97974
rect 4476 96458 4532 96460
rect 4476 96406 4478 96458
rect 4478 96406 4530 96458
rect 4530 96406 4532 96458
rect 4476 96404 4532 96406
rect 4580 96458 4636 96460
rect 4580 96406 4582 96458
rect 4582 96406 4634 96458
rect 4634 96406 4636 96458
rect 4580 96404 4636 96406
rect 4684 96458 4740 96460
rect 4684 96406 4686 96458
rect 4686 96406 4738 96458
rect 4738 96406 4740 96458
rect 4684 96404 4740 96406
rect 4476 94890 4532 94892
rect 4476 94838 4478 94890
rect 4478 94838 4530 94890
rect 4530 94838 4532 94890
rect 4476 94836 4532 94838
rect 4580 94890 4636 94892
rect 4580 94838 4582 94890
rect 4582 94838 4634 94890
rect 4634 94838 4636 94890
rect 4580 94836 4636 94838
rect 4684 94890 4740 94892
rect 4684 94838 4686 94890
rect 4686 94838 4738 94890
rect 4738 94838 4740 94890
rect 4684 94836 4740 94838
rect 4476 93322 4532 93324
rect 4476 93270 4478 93322
rect 4478 93270 4530 93322
rect 4530 93270 4532 93322
rect 4476 93268 4532 93270
rect 4580 93322 4636 93324
rect 4580 93270 4582 93322
rect 4582 93270 4634 93322
rect 4634 93270 4636 93322
rect 4580 93268 4636 93270
rect 4684 93322 4740 93324
rect 4684 93270 4686 93322
rect 4686 93270 4738 93322
rect 4738 93270 4740 93322
rect 4684 93268 4740 93270
rect 4476 91754 4532 91756
rect 4476 91702 4478 91754
rect 4478 91702 4530 91754
rect 4530 91702 4532 91754
rect 4476 91700 4532 91702
rect 4580 91754 4636 91756
rect 4580 91702 4582 91754
rect 4582 91702 4634 91754
rect 4634 91702 4636 91754
rect 4580 91700 4636 91702
rect 4684 91754 4740 91756
rect 4684 91702 4686 91754
rect 4686 91702 4738 91754
rect 4738 91702 4740 91754
rect 4684 91700 4740 91702
rect 4476 90186 4532 90188
rect 4476 90134 4478 90186
rect 4478 90134 4530 90186
rect 4530 90134 4532 90186
rect 4476 90132 4532 90134
rect 4580 90186 4636 90188
rect 4580 90134 4582 90186
rect 4582 90134 4634 90186
rect 4634 90134 4636 90186
rect 4580 90132 4636 90134
rect 4684 90186 4740 90188
rect 4684 90134 4686 90186
rect 4686 90134 4738 90186
rect 4738 90134 4740 90186
rect 4684 90132 4740 90134
rect 4476 88618 4532 88620
rect 4476 88566 4478 88618
rect 4478 88566 4530 88618
rect 4530 88566 4532 88618
rect 4476 88564 4532 88566
rect 4580 88618 4636 88620
rect 4580 88566 4582 88618
rect 4582 88566 4634 88618
rect 4634 88566 4636 88618
rect 4580 88564 4636 88566
rect 4684 88618 4740 88620
rect 4684 88566 4686 88618
rect 4686 88566 4738 88618
rect 4738 88566 4740 88618
rect 4684 88564 4740 88566
rect 4476 87050 4532 87052
rect 4476 86998 4478 87050
rect 4478 86998 4530 87050
rect 4530 86998 4532 87050
rect 4476 86996 4532 86998
rect 4580 87050 4636 87052
rect 4580 86998 4582 87050
rect 4582 86998 4634 87050
rect 4634 86998 4636 87050
rect 4580 86996 4636 86998
rect 4684 87050 4740 87052
rect 4684 86998 4686 87050
rect 4686 86998 4738 87050
rect 4738 86998 4740 87050
rect 4684 86996 4740 86998
rect 4476 85482 4532 85484
rect 4476 85430 4478 85482
rect 4478 85430 4530 85482
rect 4530 85430 4532 85482
rect 4476 85428 4532 85430
rect 4580 85482 4636 85484
rect 4580 85430 4582 85482
rect 4582 85430 4634 85482
rect 4634 85430 4636 85482
rect 4580 85428 4636 85430
rect 4684 85482 4740 85484
rect 4684 85430 4686 85482
rect 4686 85430 4738 85482
rect 4738 85430 4740 85482
rect 4684 85428 4740 85430
rect 4476 83914 4532 83916
rect 4476 83862 4478 83914
rect 4478 83862 4530 83914
rect 4530 83862 4532 83914
rect 4476 83860 4532 83862
rect 4580 83914 4636 83916
rect 4580 83862 4582 83914
rect 4582 83862 4634 83914
rect 4634 83862 4636 83914
rect 4580 83860 4636 83862
rect 4684 83914 4740 83916
rect 4684 83862 4686 83914
rect 4686 83862 4738 83914
rect 4738 83862 4740 83914
rect 4684 83860 4740 83862
rect 4476 82346 4532 82348
rect 4476 82294 4478 82346
rect 4478 82294 4530 82346
rect 4530 82294 4532 82346
rect 4476 82292 4532 82294
rect 4580 82346 4636 82348
rect 4580 82294 4582 82346
rect 4582 82294 4634 82346
rect 4634 82294 4636 82346
rect 4580 82292 4636 82294
rect 4684 82346 4740 82348
rect 4684 82294 4686 82346
rect 4686 82294 4738 82346
rect 4738 82294 4740 82346
rect 4684 82292 4740 82294
rect 4476 80778 4532 80780
rect 4476 80726 4478 80778
rect 4478 80726 4530 80778
rect 4530 80726 4532 80778
rect 4476 80724 4532 80726
rect 4580 80778 4636 80780
rect 4580 80726 4582 80778
rect 4582 80726 4634 80778
rect 4634 80726 4636 80778
rect 4580 80724 4636 80726
rect 4684 80778 4740 80780
rect 4684 80726 4686 80778
rect 4686 80726 4738 80778
rect 4738 80726 4740 80778
rect 4684 80724 4740 80726
rect 4476 79210 4532 79212
rect 4476 79158 4478 79210
rect 4478 79158 4530 79210
rect 4530 79158 4532 79210
rect 4476 79156 4532 79158
rect 4580 79210 4636 79212
rect 4580 79158 4582 79210
rect 4582 79158 4634 79210
rect 4634 79158 4636 79210
rect 4580 79156 4636 79158
rect 4684 79210 4740 79212
rect 4684 79158 4686 79210
rect 4686 79158 4738 79210
rect 4738 79158 4740 79210
rect 4684 79156 4740 79158
rect 4476 77642 4532 77644
rect 4476 77590 4478 77642
rect 4478 77590 4530 77642
rect 4530 77590 4532 77642
rect 4476 77588 4532 77590
rect 4580 77642 4636 77644
rect 4580 77590 4582 77642
rect 4582 77590 4634 77642
rect 4634 77590 4636 77642
rect 4580 77588 4636 77590
rect 4684 77642 4740 77644
rect 4684 77590 4686 77642
rect 4686 77590 4738 77642
rect 4738 77590 4740 77642
rect 4684 77588 4740 77590
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 13244 115836 13300 115892
rect 8988 20188 9044 20244
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 5964 8428 6020 8484
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 5852 3442 5908 3444
rect 5852 3390 5854 3442
rect 5854 3390 5906 3442
rect 5906 3390 5908 3442
rect 5852 3388 5908 3390
rect 8204 5852 8260 5908
rect 7868 5068 7924 5124
rect 6860 4060 6916 4116
rect 6524 3388 6580 3444
rect 8652 5906 8708 5908
rect 8652 5854 8654 5906
rect 8654 5854 8706 5906
rect 8706 5854 8708 5906
rect 8652 5852 8708 5854
rect 12572 19292 12628 19348
rect 15148 16828 15204 16884
rect 11564 6076 11620 6132
rect 8652 5122 8708 5124
rect 8652 5070 8654 5122
rect 8654 5070 8706 5122
rect 8706 5070 8708 5122
rect 8652 5068 8708 5070
rect 10668 5516 10724 5572
rect 9100 4226 9156 4228
rect 9100 4174 9102 4226
rect 9102 4174 9154 4226
rect 9154 4174 9156 4226
rect 9100 4172 9156 4174
rect 8540 4060 8596 4116
rect 9884 5010 9940 5012
rect 9884 4958 9886 5010
rect 9886 4958 9938 5010
rect 9938 4958 9940 5010
rect 9884 4956 9940 4958
rect 10444 4562 10500 4564
rect 10444 4510 10446 4562
rect 10446 4510 10498 4562
rect 10498 4510 10500 4562
rect 10444 4508 10500 4510
rect 8316 924 8372 980
rect 9884 4172 9940 4228
rect 11228 5516 11284 5572
rect 13468 6018 13524 6020
rect 13468 5966 13470 6018
rect 13470 5966 13522 6018
rect 13522 5966 13524 6018
rect 13468 5964 13524 5966
rect 11676 5068 11732 5124
rect 11452 3724 11508 3780
rect 11228 3388 11284 3444
rect 12012 5122 12068 5124
rect 12012 5070 12014 5122
rect 12014 5070 12066 5122
rect 12066 5070 12068 5122
rect 12012 5068 12068 5070
rect 12908 5068 12964 5124
rect 12124 3612 12180 3668
rect 11788 3388 11844 3444
rect 12124 3388 12180 3444
rect 11676 2604 11732 2660
rect 13692 5234 13748 5236
rect 13692 5182 13694 5234
rect 13694 5182 13746 5234
rect 13746 5182 13748 5234
rect 13692 5180 13748 5182
rect 14028 4956 14084 5012
rect 14364 5852 14420 5908
rect 14588 5346 14644 5348
rect 14588 5294 14590 5346
rect 14590 5294 14642 5346
rect 14642 5294 14644 5346
rect 14588 5292 14644 5294
rect 14252 5122 14308 5124
rect 14252 5070 14254 5122
rect 14254 5070 14306 5122
rect 14306 5070 14308 5122
rect 14252 5068 14308 5070
rect 13804 3666 13860 3668
rect 13804 3614 13806 3666
rect 13806 3614 13858 3666
rect 13858 3614 13860 3666
rect 13804 3612 13860 3614
rect 14252 3554 14308 3556
rect 14252 3502 14254 3554
rect 14254 3502 14306 3554
rect 14306 3502 14308 3554
rect 14252 3500 14308 3502
rect 14924 6466 14980 6468
rect 14924 6414 14926 6466
rect 14926 6414 14978 6466
rect 14978 6414 14980 6466
rect 14924 6412 14980 6414
rect 14812 6188 14868 6244
rect 26460 117180 26516 117236
rect 27356 117180 27412 117236
rect 28028 116508 28084 116564
rect 29484 116562 29540 116564
rect 29484 116510 29486 116562
rect 29486 116510 29538 116562
rect 29538 116510 29540 116562
rect 29484 116508 29540 116510
rect 17052 115836 17108 115892
rect 18060 116396 18116 116452
rect 16044 115666 16100 115668
rect 16044 115614 16046 115666
rect 16046 115614 16098 115666
rect 16098 115614 16100 115666
rect 16044 115612 16100 115614
rect 16716 115666 16772 115668
rect 16716 115614 16718 115666
rect 16718 115614 16770 115666
rect 16770 115614 16772 115666
rect 16716 115612 16772 115614
rect 19852 116450 19908 116452
rect 19852 116398 19854 116450
rect 19854 116398 19906 116450
rect 19906 116398 19908 116450
rect 19852 116396 19908 116398
rect 20524 116450 20580 116452
rect 20524 116398 20526 116450
rect 20526 116398 20578 116450
rect 20578 116398 20580 116450
rect 20524 116396 20580 116398
rect 19836 116058 19892 116060
rect 19836 116006 19838 116058
rect 19838 116006 19890 116058
rect 19890 116006 19892 116058
rect 19836 116004 19892 116006
rect 19940 116058 19996 116060
rect 19940 116006 19942 116058
rect 19942 116006 19994 116058
rect 19994 116006 19996 116058
rect 19940 116004 19996 116006
rect 20044 116058 20100 116060
rect 20044 116006 20046 116058
rect 20046 116006 20098 116058
rect 20098 116006 20100 116058
rect 20044 116004 20100 116006
rect 18620 115836 18676 115892
rect 20860 115666 20916 115668
rect 20860 115614 20862 115666
rect 20862 115614 20914 115666
rect 20914 115614 20916 115666
rect 20860 115612 20916 115614
rect 21532 115666 21588 115668
rect 21532 115614 21534 115666
rect 21534 115614 21586 115666
rect 21586 115614 21588 115666
rect 21532 115612 21588 115614
rect 19836 114490 19892 114492
rect 19836 114438 19838 114490
rect 19838 114438 19890 114490
rect 19890 114438 19892 114490
rect 19836 114436 19892 114438
rect 19940 114490 19996 114492
rect 19940 114438 19942 114490
rect 19942 114438 19994 114490
rect 19994 114438 19996 114490
rect 19940 114436 19996 114438
rect 20044 114490 20100 114492
rect 20044 114438 20046 114490
rect 20046 114438 20098 114490
rect 20098 114438 20100 114490
rect 20044 114436 20100 114438
rect 19836 112922 19892 112924
rect 19836 112870 19838 112922
rect 19838 112870 19890 112922
rect 19890 112870 19892 112922
rect 19836 112868 19892 112870
rect 19940 112922 19996 112924
rect 19940 112870 19942 112922
rect 19942 112870 19994 112922
rect 19994 112870 19996 112922
rect 19940 112868 19996 112870
rect 20044 112922 20100 112924
rect 20044 112870 20046 112922
rect 20046 112870 20098 112922
rect 20098 112870 20100 112922
rect 20044 112868 20100 112870
rect 19836 111354 19892 111356
rect 19836 111302 19838 111354
rect 19838 111302 19890 111354
rect 19890 111302 19892 111354
rect 19836 111300 19892 111302
rect 19940 111354 19996 111356
rect 19940 111302 19942 111354
rect 19942 111302 19994 111354
rect 19994 111302 19996 111354
rect 19940 111300 19996 111302
rect 20044 111354 20100 111356
rect 20044 111302 20046 111354
rect 20046 111302 20098 111354
rect 20098 111302 20100 111354
rect 20044 111300 20100 111302
rect 19836 109786 19892 109788
rect 19836 109734 19838 109786
rect 19838 109734 19890 109786
rect 19890 109734 19892 109786
rect 19836 109732 19892 109734
rect 19940 109786 19996 109788
rect 19940 109734 19942 109786
rect 19942 109734 19994 109786
rect 19994 109734 19996 109786
rect 19940 109732 19996 109734
rect 20044 109786 20100 109788
rect 20044 109734 20046 109786
rect 20046 109734 20098 109786
rect 20098 109734 20100 109786
rect 20044 109732 20100 109734
rect 19836 108218 19892 108220
rect 19836 108166 19838 108218
rect 19838 108166 19890 108218
rect 19890 108166 19892 108218
rect 19836 108164 19892 108166
rect 19940 108218 19996 108220
rect 19940 108166 19942 108218
rect 19942 108166 19994 108218
rect 19994 108166 19996 108218
rect 19940 108164 19996 108166
rect 20044 108218 20100 108220
rect 20044 108166 20046 108218
rect 20046 108166 20098 108218
rect 20098 108166 20100 108218
rect 20044 108164 20100 108166
rect 19836 106650 19892 106652
rect 19836 106598 19838 106650
rect 19838 106598 19890 106650
rect 19890 106598 19892 106650
rect 19836 106596 19892 106598
rect 19940 106650 19996 106652
rect 19940 106598 19942 106650
rect 19942 106598 19994 106650
rect 19994 106598 19996 106650
rect 19940 106596 19996 106598
rect 20044 106650 20100 106652
rect 20044 106598 20046 106650
rect 20046 106598 20098 106650
rect 20098 106598 20100 106650
rect 20044 106596 20100 106598
rect 19836 105082 19892 105084
rect 19836 105030 19838 105082
rect 19838 105030 19890 105082
rect 19890 105030 19892 105082
rect 19836 105028 19892 105030
rect 19940 105082 19996 105084
rect 19940 105030 19942 105082
rect 19942 105030 19994 105082
rect 19994 105030 19996 105082
rect 19940 105028 19996 105030
rect 20044 105082 20100 105084
rect 20044 105030 20046 105082
rect 20046 105030 20098 105082
rect 20098 105030 20100 105082
rect 20044 105028 20100 105030
rect 19836 103514 19892 103516
rect 19836 103462 19838 103514
rect 19838 103462 19890 103514
rect 19890 103462 19892 103514
rect 19836 103460 19892 103462
rect 19940 103514 19996 103516
rect 19940 103462 19942 103514
rect 19942 103462 19994 103514
rect 19994 103462 19996 103514
rect 19940 103460 19996 103462
rect 20044 103514 20100 103516
rect 20044 103462 20046 103514
rect 20046 103462 20098 103514
rect 20098 103462 20100 103514
rect 20044 103460 20100 103462
rect 19836 101946 19892 101948
rect 19836 101894 19838 101946
rect 19838 101894 19890 101946
rect 19890 101894 19892 101946
rect 19836 101892 19892 101894
rect 19940 101946 19996 101948
rect 19940 101894 19942 101946
rect 19942 101894 19994 101946
rect 19994 101894 19996 101946
rect 19940 101892 19996 101894
rect 20044 101946 20100 101948
rect 20044 101894 20046 101946
rect 20046 101894 20098 101946
rect 20098 101894 20100 101946
rect 20044 101892 20100 101894
rect 19836 100378 19892 100380
rect 19836 100326 19838 100378
rect 19838 100326 19890 100378
rect 19890 100326 19892 100378
rect 19836 100324 19892 100326
rect 19940 100378 19996 100380
rect 19940 100326 19942 100378
rect 19942 100326 19994 100378
rect 19994 100326 19996 100378
rect 19940 100324 19996 100326
rect 20044 100378 20100 100380
rect 20044 100326 20046 100378
rect 20046 100326 20098 100378
rect 20098 100326 20100 100378
rect 20044 100324 20100 100326
rect 19836 98810 19892 98812
rect 19836 98758 19838 98810
rect 19838 98758 19890 98810
rect 19890 98758 19892 98810
rect 19836 98756 19892 98758
rect 19940 98810 19996 98812
rect 19940 98758 19942 98810
rect 19942 98758 19994 98810
rect 19994 98758 19996 98810
rect 19940 98756 19996 98758
rect 20044 98810 20100 98812
rect 20044 98758 20046 98810
rect 20046 98758 20098 98810
rect 20098 98758 20100 98810
rect 20044 98756 20100 98758
rect 19836 97242 19892 97244
rect 19836 97190 19838 97242
rect 19838 97190 19890 97242
rect 19890 97190 19892 97242
rect 19836 97188 19892 97190
rect 19940 97242 19996 97244
rect 19940 97190 19942 97242
rect 19942 97190 19994 97242
rect 19994 97190 19996 97242
rect 19940 97188 19996 97190
rect 20044 97242 20100 97244
rect 20044 97190 20046 97242
rect 20046 97190 20098 97242
rect 20098 97190 20100 97242
rect 20044 97188 20100 97190
rect 19836 95674 19892 95676
rect 19836 95622 19838 95674
rect 19838 95622 19890 95674
rect 19890 95622 19892 95674
rect 19836 95620 19892 95622
rect 19940 95674 19996 95676
rect 19940 95622 19942 95674
rect 19942 95622 19994 95674
rect 19994 95622 19996 95674
rect 19940 95620 19996 95622
rect 20044 95674 20100 95676
rect 20044 95622 20046 95674
rect 20046 95622 20098 95674
rect 20098 95622 20100 95674
rect 20044 95620 20100 95622
rect 19836 94106 19892 94108
rect 19836 94054 19838 94106
rect 19838 94054 19890 94106
rect 19890 94054 19892 94106
rect 19836 94052 19892 94054
rect 19940 94106 19996 94108
rect 19940 94054 19942 94106
rect 19942 94054 19994 94106
rect 19994 94054 19996 94106
rect 19940 94052 19996 94054
rect 20044 94106 20100 94108
rect 20044 94054 20046 94106
rect 20046 94054 20098 94106
rect 20098 94054 20100 94106
rect 20044 94052 20100 94054
rect 19836 92538 19892 92540
rect 19836 92486 19838 92538
rect 19838 92486 19890 92538
rect 19890 92486 19892 92538
rect 19836 92484 19892 92486
rect 19940 92538 19996 92540
rect 19940 92486 19942 92538
rect 19942 92486 19994 92538
rect 19994 92486 19996 92538
rect 19940 92484 19996 92486
rect 20044 92538 20100 92540
rect 20044 92486 20046 92538
rect 20046 92486 20098 92538
rect 20098 92486 20100 92538
rect 20044 92484 20100 92486
rect 19836 90970 19892 90972
rect 19836 90918 19838 90970
rect 19838 90918 19890 90970
rect 19890 90918 19892 90970
rect 19836 90916 19892 90918
rect 19940 90970 19996 90972
rect 19940 90918 19942 90970
rect 19942 90918 19994 90970
rect 19994 90918 19996 90970
rect 19940 90916 19996 90918
rect 20044 90970 20100 90972
rect 20044 90918 20046 90970
rect 20046 90918 20098 90970
rect 20098 90918 20100 90970
rect 20044 90916 20100 90918
rect 19836 89402 19892 89404
rect 19836 89350 19838 89402
rect 19838 89350 19890 89402
rect 19890 89350 19892 89402
rect 19836 89348 19892 89350
rect 19940 89402 19996 89404
rect 19940 89350 19942 89402
rect 19942 89350 19994 89402
rect 19994 89350 19996 89402
rect 19940 89348 19996 89350
rect 20044 89402 20100 89404
rect 20044 89350 20046 89402
rect 20046 89350 20098 89402
rect 20098 89350 20100 89402
rect 20044 89348 20100 89350
rect 19836 87834 19892 87836
rect 19836 87782 19838 87834
rect 19838 87782 19890 87834
rect 19890 87782 19892 87834
rect 19836 87780 19892 87782
rect 19940 87834 19996 87836
rect 19940 87782 19942 87834
rect 19942 87782 19994 87834
rect 19994 87782 19996 87834
rect 19940 87780 19996 87782
rect 20044 87834 20100 87836
rect 20044 87782 20046 87834
rect 20046 87782 20098 87834
rect 20098 87782 20100 87834
rect 20044 87780 20100 87782
rect 19836 86266 19892 86268
rect 19836 86214 19838 86266
rect 19838 86214 19890 86266
rect 19890 86214 19892 86266
rect 19836 86212 19892 86214
rect 19940 86266 19996 86268
rect 19940 86214 19942 86266
rect 19942 86214 19994 86266
rect 19994 86214 19996 86266
rect 19940 86212 19996 86214
rect 20044 86266 20100 86268
rect 20044 86214 20046 86266
rect 20046 86214 20098 86266
rect 20098 86214 20100 86266
rect 20044 86212 20100 86214
rect 19836 84698 19892 84700
rect 19836 84646 19838 84698
rect 19838 84646 19890 84698
rect 19890 84646 19892 84698
rect 19836 84644 19892 84646
rect 19940 84698 19996 84700
rect 19940 84646 19942 84698
rect 19942 84646 19994 84698
rect 19994 84646 19996 84698
rect 19940 84644 19996 84646
rect 20044 84698 20100 84700
rect 20044 84646 20046 84698
rect 20046 84646 20098 84698
rect 20098 84646 20100 84698
rect 20044 84644 20100 84646
rect 19836 83130 19892 83132
rect 19836 83078 19838 83130
rect 19838 83078 19890 83130
rect 19890 83078 19892 83130
rect 19836 83076 19892 83078
rect 19940 83130 19996 83132
rect 19940 83078 19942 83130
rect 19942 83078 19994 83130
rect 19994 83078 19996 83130
rect 19940 83076 19996 83078
rect 20044 83130 20100 83132
rect 20044 83078 20046 83130
rect 20046 83078 20098 83130
rect 20098 83078 20100 83130
rect 20044 83076 20100 83078
rect 19836 81562 19892 81564
rect 19836 81510 19838 81562
rect 19838 81510 19890 81562
rect 19890 81510 19892 81562
rect 19836 81508 19892 81510
rect 19940 81562 19996 81564
rect 19940 81510 19942 81562
rect 19942 81510 19994 81562
rect 19994 81510 19996 81562
rect 19940 81508 19996 81510
rect 20044 81562 20100 81564
rect 20044 81510 20046 81562
rect 20046 81510 20098 81562
rect 20098 81510 20100 81562
rect 20044 81508 20100 81510
rect 19836 79994 19892 79996
rect 19836 79942 19838 79994
rect 19838 79942 19890 79994
rect 19890 79942 19892 79994
rect 19836 79940 19892 79942
rect 19940 79994 19996 79996
rect 19940 79942 19942 79994
rect 19942 79942 19994 79994
rect 19994 79942 19996 79994
rect 19940 79940 19996 79942
rect 20044 79994 20100 79996
rect 20044 79942 20046 79994
rect 20046 79942 20098 79994
rect 20098 79942 20100 79994
rect 20044 79940 20100 79942
rect 19836 78426 19892 78428
rect 19836 78374 19838 78426
rect 19838 78374 19890 78426
rect 19890 78374 19892 78426
rect 19836 78372 19892 78374
rect 19940 78426 19996 78428
rect 19940 78374 19942 78426
rect 19942 78374 19994 78426
rect 19994 78374 19996 78426
rect 19940 78372 19996 78374
rect 20044 78426 20100 78428
rect 20044 78374 20046 78426
rect 20046 78374 20098 78426
rect 20098 78374 20100 78426
rect 20044 78372 20100 78374
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 15820 8652 15876 8708
rect 14924 6018 14980 6020
rect 14924 5966 14926 6018
rect 14926 5966 14978 6018
rect 14978 5966 14980 6018
rect 14924 5964 14980 5966
rect 14812 5180 14868 5236
rect 15036 5180 15092 5236
rect 16828 18508 16884 18564
rect 14700 3500 14756 3556
rect 14812 3388 14868 3444
rect 14588 3330 14644 3332
rect 14588 3278 14590 3330
rect 14590 3278 14642 3330
rect 14642 3278 14644 3330
rect 14588 3276 14644 3278
rect 15820 5292 15876 5348
rect 16380 6300 16436 6356
rect 16604 5906 16660 5908
rect 16604 5854 16606 5906
rect 16606 5854 16658 5906
rect 16658 5854 16660 5906
rect 16604 5852 16660 5854
rect 16044 5292 16100 5348
rect 17388 6300 17444 6356
rect 17724 6188 17780 6244
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 23100 18620 23156 18676
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21980 13580 22036 13636
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 18620 10108 18676 10164
rect 18284 7308 18340 7364
rect 17388 5852 17444 5908
rect 17164 4396 17220 4452
rect 16156 4172 16212 4228
rect 18396 6188 18452 6244
rect 18396 6018 18452 6020
rect 18396 5966 18398 6018
rect 18398 5966 18450 6018
rect 18450 5966 18452 6018
rect 18396 5964 18452 5966
rect 17836 4226 17892 4228
rect 17836 4174 17838 4226
rect 17838 4174 17890 4226
rect 17890 4174 17892 4226
rect 17836 4172 17892 4174
rect 15820 3948 15876 4004
rect 17724 3948 17780 4004
rect 16604 3500 16660 3556
rect 16044 3442 16100 3444
rect 16044 3390 16046 3442
rect 16046 3390 16098 3442
rect 16098 3390 16100 3442
rect 16044 3388 16100 3390
rect 17164 3388 17220 3444
rect 17836 3442 17892 3444
rect 17836 3390 17838 3442
rect 17838 3390 17890 3442
rect 17890 3390 17892 3442
rect 17836 3388 17892 3390
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19292 7308 19348 7364
rect 18844 6300 18900 6356
rect 18732 5292 18788 5348
rect 18396 4396 18452 4452
rect 19068 5180 19124 5236
rect 19180 6300 19236 6356
rect 19180 4844 19236 4900
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19964 6914 20020 6916
rect 19964 6862 19966 6914
rect 19966 6862 20018 6914
rect 20018 6862 20020 6914
rect 19964 6860 20020 6862
rect 20188 6524 20244 6580
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20636 6524 20692 6580
rect 21532 7362 21588 7364
rect 21532 7310 21534 7362
rect 21534 7310 21586 7362
rect 21586 7310 21588 7362
rect 21532 7308 21588 7310
rect 22764 9324 22820 9380
rect 22428 7362 22484 7364
rect 22428 7310 22430 7362
rect 22430 7310 22482 7362
rect 22482 7310 22484 7362
rect 22428 7308 22484 7310
rect 21980 7196 22036 7252
rect 21980 6860 22036 6916
rect 22092 7084 22148 7140
rect 21532 6578 21588 6580
rect 21532 6526 21534 6578
rect 21534 6526 21586 6578
rect 21586 6526 21588 6578
rect 21532 6524 21588 6526
rect 20076 5964 20132 6020
rect 19852 5794 19908 5796
rect 19852 5742 19854 5794
rect 19854 5742 19906 5794
rect 19906 5742 19908 5794
rect 19852 5740 19908 5742
rect 19292 3612 19348 3668
rect 18172 2716 18228 2772
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20524 5740 20580 5796
rect 19740 3442 19796 3444
rect 19740 3390 19742 3442
rect 19742 3390 19794 3442
rect 19794 3390 19796 3442
rect 19740 3388 19796 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21196 5740 21252 5796
rect 21644 5180 21700 5236
rect 20636 3554 20692 3556
rect 20636 3502 20638 3554
rect 20638 3502 20690 3554
rect 20690 3502 20692 3554
rect 20636 3500 20692 3502
rect 21084 3388 21140 3444
rect 21644 1596 21700 1652
rect 21868 5234 21924 5236
rect 21868 5182 21870 5234
rect 21870 5182 21922 5234
rect 21922 5182 21924 5234
rect 21868 5180 21924 5182
rect 22540 6524 22596 6580
rect 21980 3500 22036 3556
rect 21756 1148 21812 1204
rect 22428 3500 22484 3556
rect 22876 6524 22932 6580
rect 24444 12796 24500 12852
rect 23212 6300 23268 6356
rect 22876 4338 22932 4340
rect 22876 4286 22878 4338
rect 22878 4286 22930 4338
rect 22930 4286 22932 4338
rect 22876 4284 22932 4286
rect 23548 6300 23604 6356
rect 24220 7084 24276 7140
rect 24332 7196 24388 7252
rect 31164 116620 31220 116676
rect 31948 116620 32004 116676
rect 35196 116842 35252 116844
rect 35196 116790 35198 116842
rect 35198 116790 35250 116842
rect 35250 116790 35252 116842
rect 35196 116788 35252 116790
rect 35300 116842 35356 116844
rect 35300 116790 35302 116842
rect 35302 116790 35354 116842
rect 35354 116790 35356 116842
rect 35300 116788 35356 116790
rect 35404 116842 35460 116844
rect 35404 116790 35406 116842
rect 35406 116790 35458 116842
rect 35458 116790 35460 116842
rect 35404 116788 35460 116790
rect 32732 116508 32788 116564
rect 33628 116562 33684 116564
rect 33628 116510 33630 116562
rect 33630 116510 33682 116562
rect 33682 116510 33684 116562
rect 33628 116508 33684 116510
rect 25564 115666 25620 115668
rect 25564 115614 25566 115666
rect 25566 115614 25618 115666
rect 25618 115614 25620 115666
rect 25564 115612 25620 115614
rect 26236 115666 26292 115668
rect 26236 115614 26238 115666
rect 26238 115614 26290 115666
rect 26290 115614 26292 115666
rect 26236 115612 26292 115614
rect 30268 115666 30324 115668
rect 30268 115614 30270 115666
rect 30270 115614 30322 115666
rect 30322 115614 30324 115666
rect 30268 115612 30324 115614
rect 30940 115666 30996 115668
rect 30940 115614 30942 115666
rect 30942 115614 30994 115666
rect 30994 115614 30996 115666
rect 30940 115612 30996 115614
rect 25788 22540 25844 22596
rect 34636 115666 34692 115668
rect 34636 115614 34638 115666
rect 34638 115614 34690 115666
rect 34690 115614 34692 115666
rect 34636 115612 34692 115614
rect 33628 22428 33684 22484
rect 26908 16716 26964 16772
rect 24892 6130 24948 6132
rect 24892 6078 24894 6130
rect 24894 6078 24946 6130
rect 24946 6078 24948 6130
rect 24892 6076 24948 6078
rect 23772 5180 23828 5236
rect 23436 4396 23492 4452
rect 23324 4284 23380 4340
rect 23660 3442 23716 3444
rect 23660 3390 23662 3442
rect 23662 3390 23714 3442
rect 23714 3390 23716 3442
rect 23660 3388 23716 3390
rect 24108 3500 24164 3556
rect 24556 3554 24612 3556
rect 24556 3502 24558 3554
rect 24558 3502 24610 3554
rect 24610 3502 24612 3554
rect 24556 3500 24612 3502
rect 25340 4284 25396 4340
rect 25452 3724 25508 3780
rect 26796 7756 26852 7812
rect 25676 7308 25732 7364
rect 25676 6076 25732 6132
rect 29708 16044 29764 16100
rect 28476 13692 28532 13748
rect 27804 8316 27860 8372
rect 27804 7756 27860 7812
rect 27804 6802 27860 6804
rect 27804 6750 27806 6802
rect 27806 6750 27858 6802
rect 27858 6750 27860 6802
rect 27804 6748 27860 6750
rect 26908 6076 26964 6132
rect 27580 4450 27636 4452
rect 27580 4398 27582 4450
rect 27582 4398 27634 4450
rect 27634 4398 27636 4450
rect 27580 4396 27636 4398
rect 27132 3724 27188 3780
rect 26124 3388 26180 3444
rect 24780 1036 24836 1092
rect 27244 3500 27300 3556
rect 27468 3388 27524 3444
rect 28252 3554 28308 3556
rect 28252 3502 28254 3554
rect 28254 3502 28306 3554
rect 28306 3502 28308 3554
rect 28252 3500 28308 3502
rect 28140 3388 28196 3444
rect 29148 7644 29204 7700
rect 29036 6076 29092 6132
rect 29148 6748 29204 6804
rect 28588 4396 28644 4452
rect 28588 4226 28644 4228
rect 28588 4174 28590 4226
rect 28590 4174 28642 4226
rect 28642 4174 28644 4226
rect 28588 4172 28644 4174
rect 29148 4172 29204 4228
rect 29260 3500 29316 3556
rect 29484 3724 29540 3780
rect 29932 12124 29988 12180
rect 30716 9548 30772 9604
rect 30604 6636 30660 6692
rect 30044 3724 30100 3780
rect 30604 6076 30660 6132
rect 31052 7308 31108 7364
rect 30940 6412 30996 6468
rect 32956 17612 33012 17668
rect 32844 9548 32900 9604
rect 32172 9042 32228 9044
rect 32172 8990 32174 9042
rect 32174 8990 32226 9042
rect 32226 8990 32228 9042
rect 32172 8988 32228 8990
rect 32284 7586 32340 7588
rect 32284 7534 32286 7586
rect 32286 7534 32338 7586
rect 32338 7534 32340 7586
rect 32284 7532 32340 7534
rect 31276 7084 31332 7140
rect 31052 6188 31108 6244
rect 32844 7196 32900 7252
rect 31500 5852 31556 5908
rect 31612 5794 31668 5796
rect 31612 5742 31614 5794
rect 31614 5742 31666 5794
rect 31666 5742 31668 5794
rect 31612 5740 31668 5742
rect 30492 3388 30548 3444
rect 30604 3500 30660 3556
rect 30940 3442 30996 3444
rect 30940 3390 30942 3442
rect 30942 3390 30994 3442
rect 30994 3390 30996 3442
rect 30940 3388 30996 3390
rect 30828 1260 30884 1316
rect 32060 6412 32116 6468
rect 38892 116284 38948 116340
rect 39340 116338 39396 116340
rect 39340 116286 39342 116338
rect 39342 116286 39394 116338
rect 39394 116286 39396 116338
rect 39340 116284 39396 116286
rect 49980 117180 50036 117236
rect 50876 117180 50932 117236
rect 54684 116956 54740 117012
rect 55468 116956 55524 117012
rect 51548 116508 51604 116564
rect 53004 116562 53060 116564
rect 53004 116510 53006 116562
rect 53006 116510 53058 116562
rect 53058 116510 53060 116562
rect 53004 116508 53060 116510
rect 56252 116508 56308 116564
rect 57148 116562 57204 116564
rect 57148 116510 57150 116562
rect 57150 116510 57202 116562
rect 57202 116510 57204 116562
rect 57148 116508 57204 116510
rect 35868 115836 35924 115892
rect 36764 115836 36820 115892
rect 35196 115666 35252 115668
rect 35196 115614 35198 115666
rect 35198 115614 35250 115666
rect 35250 115614 35252 115666
rect 35196 115612 35252 115614
rect 40684 115836 40740 115892
rect 42252 115836 42308 115892
rect 39676 115666 39732 115668
rect 39676 115614 39678 115666
rect 39678 115614 39730 115666
rect 39730 115614 39732 115666
rect 39676 115612 39732 115614
rect 40236 115666 40292 115668
rect 40236 115614 40238 115666
rect 40238 115614 40290 115666
rect 40290 115614 40292 115666
rect 40236 115612 40292 115614
rect 35196 115274 35252 115276
rect 35196 115222 35198 115274
rect 35198 115222 35250 115274
rect 35250 115222 35252 115274
rect 35196 115220 35252 115222
rect 35300 115274 35356 115276
rect 35300 115222 35302 115274
rect 35302 115222 35354 115274
rect 35354 115222 35356 115274
rect 35300 115220 35356 115222
rect 35404 115274 35460 115276
rect 35404 115222 35406 115274
rect 35406 115222 35458 115274
rect 35458 115222 35460 115274
rect 35404 115220 35460 115222
rect 35196 113706 35252 113708
rect 35196 113654 35198 113706
rect 35198 113654 35250 113706
rect 35250 113654 35252 113706
rect 35196 113652 35252 113654
rect 35300 113706 35356 113708
rect 35300 113654 35302 113706
rect 35302 113654 35354 113706
rect 35354 113654 35356 113706
rect 35300 113652 35356 113654
rect 35404 113706 35460 113708
rect 35404 113654 35406 113706
rect 35406 113654 35458 113706
rect 35458 113654 35460 113706
rect 35404 113652 35460 113654
rect 35196 112138 35252 112140
rect 35196 112086 35198 112138
rect 35198 112086 35250 112138
rect 35250 112086 35252 112138
rect 35196 112084 35252 112086
rect 35300 112138 35356 112140
rect 35300 112086 35302 112138
rect 35302 112086 35354 112138
rect 35354 112086 35356 112138
rect 35300 112084 35356 112086
rect 35404 112138 35460 112140
rect 35404 112086 35406 112138
rect 35406 112086 35458 112138
rect 35458 112086 35460 112138
rect 35404 112084 35460 112086
rect 35196 110570 35252 110572
rect 35196 110518 35198 110570
rect 35198 110518 35250 110570
rect 35250 110518 35252 110570
rect 35196 110516 35252 110518
rect 35300 110570 35356 110572
rect 35300 110518 35302 110570
rect 35302 110518 35354 110570
rect 35354 110518 35356 110570
rect 35300 110516 35356 110518
rect 35404 110570 35460 110572
rect 35404 110518 35406 110570
rect 35406 110518 35458 110570
rect 35458 110518 35460 110570
rect 35404 110516 35460 110518
rect 35196 109002 35252 109004
rect 35196 108950 35198 109002
rect 35198 108950 35250 109002
rect 35250 108950 35252 109002
rect 35196 108948 35252 108950
rect 35300 109002 35356 109004
rect 35300 108950 35302 109002
rect 35302 108950 35354 109002
rect 35354 108950 35356 109002
rect 35300 108948 35356 108950
rect 35404 109002 35460 109004
rect 35404 108950 35406 109002
rect 35406 108950 35458 109002
rect 35458 108950 35460 109002
rect 35404 108948 35460 108950
rect 35196 107434 35252 107436
rect 35196 107382 35198 107434
rect 35198 107382 35250 107434
rect 35250 107382 35252 107434
rect 35196 107380 35252 107382
rect 35300 107434 35356 107436
rect 35300 107382 35302 107434
rect 35302 107382 35354 107434
rect 35354 107382 35356 107434
rect 35300 107380 35356 107382
rect 35404 107434 35460 107436
rect 35404 107382 35406 107434
rect 35406 107382 35458 107434
rect 35458 107382 35460 107434
rect 35404 107380 35460 107382
rect 35196 105866 35252 105868
rect 35196 105814 35198 105866
rect 35198 105814 35250 105866
rect 35250 105814 35252 105866
rect 35196 105812 35252 105814
rect 35300 105866 35356 105868
rect 35300 105814 35302 105866
rect 35302 105814 35354 105866
rect 35354 105814 35356 105866
rect 35300 105812 35356 105814
rect 35404 105866 35460 105868
rect 35404 105814 35406 105866
rect 35406 105814 35458 105866
rect 35458 105814 35460 105866
rect 35404 105812 35460 105814
rect 35196 104298 35252 104300
rect 35196 104246 35198 104298
rect 35198 104246 35250 104298
rect 35250 104246 35252 104298
rect 35196 104244 35252 104246
rect 35300 104298 35356 104300
rect 35300 104246 35302 104298
rect 35302 104246 35354 104298
rect 35354 104246 35356 104298
rect 35300 104244 35356 104246
rect 35404 104298 35460 104300
rect 35404 104246 35406 104298
rect 35406 104246 35458 104298
rect 35458 104246 35460 104298
rect 35404 104244 35460 104246
rect 35196 102730 35252 102732
rect 35196 102678 35198 102730
rect 35198 102678 35250 102730
rect 35250 102678 35252 102730
rect 35196 102676 35252 102678
rect 35300 102730 35356 102732
rect 35300 102678 35302 102730
rect 35302 102678 35354 102730
rect 35354 102678 35356 102730
rect 35300 102676 35356 102678
rect 35404 102730 35460 102732
rect 35404 102678 35406 102730
rect 35406 102678 35458 102730
rect 35458 102678 35460 102730
rect 35404 102676 35460 102678
rect 35196 101162 35252 101164
rect 35196 101110 35198 101162
rect 35198 101110 35250 101162
rect 35250 101110 35252 101162
rect 35196 101108 35252 101110
rect 35300 101162 35356 101164
rect 35300 101110 35302 101162
rect 35302 101110 35354 101162
rect 35354 101110 35356 101162
rect 35300 101108 35356 101110
rect 35404 101162 35460 101164
rect 35404 101110 35406 101162
rect 35406 101110 35458 101162
rect 35458 101110 35460 101162
rect 35404 101108 35460 101110
rect 35196 99594 35252 99596
rect 35196 99542 35198 99594
rect 35198 99542 35250 99594
rect 35250 99542 35252 99594
rect 35196 99540 35252 99542
rect 35300 99594 35356 99596
rect 35300 99542 35302 99594
rect 35302 99542 35354 99594
rect 35354 99542 35356 99594
rect 35300 99540 35356 99542
rect 35404 99594 35460 99596
rect 35404 99542 35406 99594
rect 35406 99542 35458 99594
rect 35458 99542 35460 99594
rect 35404 99540 35460 99542
rect 35196 98026 35252 98028
rect 35196 97974 35198 98026
rect 35198 97974 35250 98026
rect 35250 97974 35252 98026
rect 35196 97972 35252 97974
rect 35300 98026 35356 98028
rect 35300 97974 35302 98026
rect 35302 97974 35354 98026
rect 35354 97974 35356 98026
rect 35300 97972 35356 97974
rect 35404 98026 35460 98028
rect 35404 97974 35406 98026
rect 35406 97974 35458 98026
rect 35458 97974 35460 98026
rect 35404 97972 35460 97974
rect 35196 96458 35252 96460
rect 35196 96406 35198 96458
rect 35198 96406 35250 96458
rect 35250 96406 35252 96458
rect 35196 96404 35252 96406
rect 35300 96458 35356 96460
rect 35300 96406 35302 96458
rect 35302 96406 35354 96458
rect 35354 96406 35356 96458
rect 35300 96404 35356 96406
rect 35404 96458 35460 96460
rect 35404 96406 35406 96458
rect 35406 96406 35458 96458
rect 35458 96406 35460 96458
rect 35404 96404 35460 96406
rect 35196 94890 35252 94892
rect 35196 94838 35198 94890
rect 35198 94838 35250 94890
rect 35250 94838 35252 94890
rect 35196 94836 35252 94838
rect 35300 94890 35356 94892
rect 35300 94838 35302 94890
rect 35302 94838 35354 94890
rect 35354 94838 35356 94890
rect 35300 94836 35356 94838
rect 35404 94890 35460 94892
rect 35404 94838 35406 94890
rect 35406 94838 35458 94890
rect 35458 94838 35460 94890
rect 35404 94836 35460 94838
rect 35196 93322 35252 93324
rect 35196 93270 35198 93322
rect 35198 93270 35250 93322
rect 35250 93270 35252 93322
rect 35196 93268 35252 93270
rect 35300 93322 35356 93324
rect 35300 93270 35302 93322
rect 35302 93270 35354 93322
rect 35354 93270 35356 93322
rect 35300 93268 35356 93270
rect 35404 93322 35460 93324
rect 35404 93270 35406 93322
rect 35406 93270 35458 93322
rect 35458 93270 35460 93322
rect 35404 93268 35460 93270
rect 35196 91754 35252 91756
rect 35196 91702 35198 91754
rect 35198 91702 35250 91754
rect 35250 91702 35252 91754
rect 35196 91700 35252 91702
rect 35300 91754 35356 91756
rect 35300 91702 35302 91754
rect 35302 91702 35354 91754
rect 35354 91702 35356 91754
rect 35300 91700 35356 91702
rect 35404 91754 35460 91756
rect 35404 91702 35406 91754
rect 35406 91702 35458 91754
rect 35458 91702 35460 91754
rect 35404 91700 35460 91702
rect 35196 90186 35252 90188
rect 35196 90134 35198 90186
rect 35198 90134 35250 90186
rect 35250 90134 35252 90186
rect 35196 90132 35252 90134
rect 35300 90186 35356 90188
rect 35300 90134 35302 90186
rect 35302 90134 35354 90186
rect 35354 90134 35356 90186
rect 35300 90132 35356 90134
rect 35404 90186 35460 90188
rect 35404 90134 35406 90186
rect 35406 90134 35458 90186
rect 35458 90134 35460 90186
rect 35404 90132 35460 90134
rect 35196 88618 35252 88620
rect 35196 88566 35198 88618
rect 35198 88566 35250 88618
rect 35250 88566 35252 88618
rect 35196 88564 35252 88566
rect 35300 88618 35356 88620
rect 35300 88566 35302 88618
rect 35302 88566 35354 88618
rect 35354 88566 35356 88618
rect 35300 88564 35356 88566
rect 35404 88618 35460 88620
rect 35404 88566 35406 88618
rect 35406 88566 35458 88618
rect 35458 88566 35460 88618
rect 35404 88564 35460 88566
rect 35196 87050 35252 87052
rect 35196 86998 35198 87050
rect 35198 86998 35250 87050
rect 35250 86998 35252 87050
rect 35196 86996 35252 86998
rect 35300 87050 35356 87052
rect 35300 86998 35302 87050
rect 35302 86998 35354 87050
rect 35354 86998 35356 87050
rect 35300 86996 35356 86998
rect 35404 87050 35460 87052
rect 35404 86998 35406 87050
rect 35406 86998 35458 87050
rect 35458 86998 35460 87050
rect 35404 86996 35460 86998
rect 35196 85482 35252 85484
rect 35196 85430 35198 85482
rect 35198 85430 35250 85482
rect 35250 85430 35252 85482
rect 35196 85428 35252 85430
rect 35300 85482 35356 85484
rect 35300 85430 35302 85482
rect 35302 85430 35354 85482
rect 35354 85430 35356 85482
rect 35300 85428 35356 85430
rect 35404 85482 35460 85484
rect 35404 85430 35406 85482
rect 35406 85430 35458 85482
rect 35458 85430 35460 85482
rect 35404 85428 35460 85430
rect 35196 83914 35252 83916
rect 35196 83862 35198 83914
rect 35198 83862 35250 83914
rect 35250 83862 35252 83914
rect 35196 83860 35252 83862
rect 35300 83914 35356 83916
rect 35300 83862 35302 83914
rect 35302 83862 35354 83914
rect 35354 83862 35356 83914
rect 35300 83860 35356 83862
rect 35404 83914 35460 83916
rect 35404 83862 35406 83914
rect 35406 83862 35458 83914
rect 35458 83862 35460 83914
rect 35404 83860 35460 83862
rect 35196 82346 35252 82348
rect 35196 82294 35198 82346
rect 35198 82294 35250 82346
rect 35250 82294 35252 82346
rect 35196 82292 35252 82294
rect 35300 82346 35356 82348
rect 35300 82294 35302 82346
rect 35302 82294 35354 82346
rect 35354 82294 35356 82346
rect 35300 82292 35356 82294
rect 35404 82346 35460 82348
rect 35404 82294 35406 82346
rect 35406 82294 35458 82346
rect 35458 82294 35460 82346
rect 35404 82292 35460 82294
rect 35196 80778 35252 80780
rect 35196 80726 35198 80778
rect 35198 80726 35250 80778
rect 35250 80726 35252 80778
rect 35196 80724 35252 80726
rect 35300 80778 35356 80780
rect 35300 80726 35302 80778
rect 35302 80726 35354 80778
rect 35354 80726 35356 80778
rect 35300 80724 35356 80726
rect 35404 80778 35460 80780
rect 35404 80726 35406 80778
rect 35406 80726 35458 80778
rect 35458 80726 35460 80778
rect 35404 80724 35460 80726
rect 35196 79210 35252 79212
rect 35196 79158 35198 79210
rect 35198 79158 35250 79210
rect 35250 79158 35252 79210
rect 35196 79156 35252 79158
rect 35300 79210 35356 79212
rect 35300 79158 35302 79210
rect 35302 79158 35354 79210
rect 35354 79158 35356 79210
rect 35300 79156 35356 79158
rect 35404 79210 35460 79212
rect 35404 79158 35406 79210
rect 35406 79158 35458 79210
rect 35458 79158 35460 79210
rect 35404 79156 35460 79158
rect 35196 77642 35252 77644
rect 35196 77590 35198 77642
rect 35198 77590 35250 77642
rect 35250 77590 35252 77642
rect 35196 77588 35252 77590
rect 35300 77642 35356 77644
rect 35300 77590 35302 77642
rect 35302 77590 35354 77642
rect 35354 77590 35356 77642
rect 35300 77588 35356 77590
rect 35404 77642 35460 77644
rect 35404 77590 35406 77642
rect 35406 77590 35458 77642
rect 35458 77590 35460 77642
rect 35404 77588 35460 77590
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 48076 116450 48132 116452
rect 48076 116398 48078 116450
rect 48078 116398 48130 116450
rect 48130 116398 48132 116450
rect 48076 116396 48132 116398
rect 48748 116396 48804 116452
rect 44380 115666 44436 115668
rect 44380 115614 44382 115666
rect 44382 115614 44434 115666
rect 44434 115614 44436 115666
rect 44380 115612 44436 115614
rect 45052 115666 45108 115668
rect 45052 115614 45054 115666
rect 45054 115614 45106 115666
rect 45106 115614 45108 115666
rect 45052 115612 45108 115614
rect 48748 115666 48804 115668
rect 48748 115614 48750 115666
rect 48750 115614 48802 115666
rect 48802 115614 48804 115666
rect 48748 115612 48804 115614
rect 50556 116058 50612 116060
rect 50556 116006 50558 116058
rect 50558 116006 50610 116058
rect 50610 116006 50612 116058
rect 50556 116004 50612 116006
rect 50660 116058 50716 116060
rect 50660 116006 50662 116058
rect 50662 116006 50714 116058
rect 50714 116006 50716 116058
rect 50660 116004 50716 116006
rect 50764 116058 50820 116060
rect 50764 116006 50766 116058
rect 50766 116006 50818 116058
rect 50818 116006 50820 116058
rect 50764 116004 50820 116006
rect 57932 116060 57988 116116
rect 58380 116060 58436 116116
rect 59388 115836 59444 115892
rect 60284 115836 60340 115892
rect 53788 115724 53844 115780
rect 49756 115666 49812 115668
rect 49756 115614 49758 115666
rect 49758 115614 49810 115666
rect 49810 115614 49812 115666
rect 49756 115612 49812 115614
rect 50556 114490 50612 114492
rect 50556 114438 50558 114490
rect 50558 114438 50610 114490
rect 50610 114438 50612 114490
rect 50556 114436 50612 114438
rect 50660 114490 50716 114492
rect 50660 114438 50662 114490
rect 50662 114438 50714 114490
rect 50714 114438 50716 114490
rect 50660 114436 50716 114438
rect 50764 114490 50820 114492
rect 50764 114438 50766 114490
rect 50766 114438 50818 114490
rect 50818 114438 50820 114490
rect 50764 114436 50820 114438
rect 50556 112922 50612 112924
rect 50556 112870 50558 112922
rect 50558 112870 50610 112922
rect 50610 112870 50612 112922
rect 50556 112868 50612 112870
rect 50660 112922 50716 112924
rect 50660 112870 50662 112922
rect 50662 112870 50714 112922
rect 50714 112870 50716 112922
rect 50660 112868 50716 112870
rect 50764 112922 50820 112924
rect 50764 112870 50766 112922
rect 50766 112870 50818 112922
rect 50818 112870 50820 112922
rect 50764 112868 50820 112870
rect 50556 111354 50612 111356
rect 50556 111302 50558 111354
rect 50558 111302 50610 111354
rect 50610 111302 50612 111354
rect 50556 111300 50612 111302
rect 50660 111354 50716 111356
rect 50660 111302 50662 111354
rect 50662 111302 50714 111354
rect 50714 111302 50716 111354
rect 50660 111300 50716 111302
rect 50764 111354 50820 111356
rect 50764 111302 50766 111354
rect 50766 111302 50818 111354
rect 50818 111302 50820 111354
rect 50764 111300 50820 111302
rect 50556 109786 50612 109788
rect 50556 109734 50558 109786
rect 50558 109734 50610 109786
rect 50610 109734 50612 109786
rect 50556 109732 50612 109734
rect 50660 109786 50716 109788
rect 50660 109734 50662 109786
rect 50662 109734 50714 109786
rect 50714 109734 50716 109786
rect 50660 109732 50716 109734
rect 50764 109786 50820 109788
rect 50764 109734 50766 109786
rect 50766 109734 50818 109786
rect 50818 109734 50820 109786
rect 50764 109732 50820 109734
rect 50556 108218 50612 108220
rect 50556 108166 50558 108218
rect 50558 108166 50610 108218
rect 50610 108166 50612 108218
rect 50556 108164 50612 108166
rect 50660 108218 50716 108220
rect 50660 108166 50662 108218
rect 50662 108166 50714 108218
rect 50714 108166 50716 108218
rect 50660 108164 50716 108166
rect 50764 108218 50820 108220
rect 50764 108166 50766 108218
rect 50766 108166 50818 108218
rect 50818 108166 50820 108218
rect 50764 108164 50820 108166
rect 50556 106650 50612 106652
rect 50556 106598 50558 106650
rect 50558 106598 50610 106650
rect 50610 106598 50612 106650
rect 50556 106596 50612 106598
rect 50660 106650 50716 106652
rect 50660 106598 50662 106650
rect 50662 106598 50714 106650
rect 50714 106598 50716 106650
rect 50660 106596 50716 106598
rect 50764 106650 50820 106652
rect 50764 106598 50766 106650
rect 50766 106598 50818 106650
rect 50818 106598 50820 106650
rect 50764 106596 50820 106598
rect 50556 105082 50612 105084
rect 50556 105030 50558 105082
rect 50558 105030 50610 105082
rect 50610 105030 50612 105082
rect 50556 105028 50612 105030
rect 50660 105082 50716 105084
rect 50660 105030 50662 105082
rect 50662 105030 50714 105082
rect 50714 105030 50716 105082
rect 50660 105028 50716 105030
rect 50764 105082 50820 105084
rect 50764 105030 50766 105082
rect 50766 105030 50818 105082
rect 50818 105030 50820 105082
rect 50764 105028 50820 105030
rect 50556 103514 50612 103516
rect 50556 103462 50558 103514
rect 50558 103462 50610 103514
rect 50610 103462 50612 103514
rect 50556 103460 50612 103462
rect 50660 103514 50716 103516
rect 50660 103462 50662 103514
rect 50662 103462 50714 103514
rect 50714 103462 50716 103514
rect 50660 103460 50716 103462
rect 50764 103514 50820 103516
rect 50764 103462 50766 103514
rect 50766 103462 50818 103514
rect 50818 103462 50820 103514
rect 50764 103460 50820 103462
rect 55132 115778 55188 115780
rect 55132 115726 55134 115778
rect 55134 115726 55186 115778
rect 55186 115726 55188 115778
rect 55132 115724 55188 115726
rect 54460 115666 54516 115668
rect 54460 115614 54462 115666
rect 54462 115614 54514 115666
rect 54514 115614 54516 115666
rect 54460 115612 54516 115614
rect 53788 115554 53844 115556
rect 53788 115502 53790 115554
rect 53790 115502 53842 115554
rect 53842 115502 53844 115554
rect 53788 115500 53844 115502
rect 58156 115554 58212 115556
rect 58156 115502 58158 115554
rect 58158 115502 58210 115554
rect 58210 115502 58212 115554
rect 58156 115500 58212 115502
rect 58716 115500 58772 115556
rect 43708 29372 43764 29428
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 45276 27244 45332 27300
rect 41020 27020 41076 27076
rect 40012 26908 40068 26964
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 38556 22988 38612 23044
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34860 22428 34916 22484
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 33628 16716 33684 16772
rect 35084 19404 35140 19460
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 37884 15372 37940 15428
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 36876 12348 36932 12404
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 33964 9602 34020 9604
rect 33964 9550 33966 9602
rect 33966 9550 34018 9602
rect 34018 9550 34020 9602
rect 33964 9548 34020 9550
rect 33516 9100 33572 9156
rect 34636 9154 34692 9156
rect 34636 9102 34638 9154
rect 34638 9102 34690 9154
rect 34690 9102 34692 9154
rect 34636 9100 34692 9102
rect 33740 9042 33796 9044
rect 33740 8990 33742 9042
rect 33742 8990 33794 9042
rect 33794 8990 33796 9042
rect 33740 8988 33796 8990
rect 34076 9042 34132 9044
rect 34076 8990 34078 9042
rect 34078 8990 34130 9042
rect 34130 8990 34132 9042
rect 34076 8988 34132 8990
rect 33068 7420 33124 7476
rect 32620 5906 32676 5908
rect 32620 5854 32622 5906
rect 32622 5854 32674 5906
rect 32674 5854 32676 5906
rect 32620 5852 32676 5854
rect 32060 5628 32116 5684
rect 33516 7474 33572 7476
rect 33516 7422 33518 7474
rect 33518 7422 33570 7474
rect 33570 7422 33572 7474
rect 33516 7420 33572 7422
rect 34188 7196 34244 7252
rect 34188 6578 34244 6580
rect 34188 6526 34190 6578
rect 34190 6526 34242 6578
rect 34242 6526 34244 6578
rect 34188 6524 34244 6526
rect 34188 6018 34244 6020
rect 34188 5966 34190 6018
rect 34190 5966 34242 6018
rect 34242 5966 34244 6018
rect 34188 5964 34244 5966
rect 33068 5516 33124 5572
rect 31724 4956 31780 5012
rect 32508 4844 32564 4900
rect 31500 3442 31556 3444
rect 31500 3390 31502 3442
rect 31502 3390 31554 3442
rect 31554 3390 31556 3442
rect 31500 3388 31556 3390
rect 32060 3388 32116 3444
rect 32284 3724 32340 3780
rect 33516 4844 33572 4900
rect 33852 4844 33908 4900
rect 33964 5852 34020 5908
rect 33516 4562 33572 4564
rect 33516 4510 33518 4562
rect 33518 4510 33570 4562
rect 33570 4510 33572 4562
rect 33516 4508 33572 4510
rect 32844 4338 32900 4340
rect 32844 4286 32846 4338
rect 32846 4286 32898 4338
rect 32898 4286 32900 4338
rect 32844 4284 32900 4286
rect 32844 3388 32900 3444
rect 33516 3442 33572 3444
rect 33516 3390 33518 3442
rect 33518 3390 33570 3442
rect 33570 3390 33572 3442
rect 33516 3388 33572 3390
rect 34524 7868 34580 7924
rect 34748 7868 34804 7924
rect 36316 9996 36372 10052
rect 35420 8988 35476 9044
rect 35084 8876 35140 8932
rect 35868 8930 35924 8932
rect 35868 8878 35870 8930
rect 35870 8878 35922 8930
rect 35922 8878 35924 8930
rect 35868 8876 35924 8878
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35084 8258 35140 8260
rect 35084 8206 35086 8258
rect 35086 8206 35138 8258
rect 35138 8206 35140 8258
rect 35084 8204 35140 8206
rect 35420 7532 35476 7588
rect 35308 7362 35364 7364
rect 35308 7310 35310 7362
rect 35310 7310 35362 7362
rect 35362 7310 35364 7362
rect 35308 7308 35364 7310
rect 36540 9714 36596 9716
rect 36540 9662 36542 9714
rect 36542 9662 36594 9714
rect 36594 9662 36596 9714
rect 36540 9660 36596 9662
rect 36092 7474 36148 7476
rect 36092 7422 36094 7474
rect 36094 7422 36146 7474
rect 36146 7422 36148 7474
rect 36092 7420 36148 7422
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34860 6690 34916 6692
rect 34860 6638 34862 6690
rect 34862 6638 34914 6690
rect 34914 6638 34916 6690
rect 34860 6636 34916 6638
rect 34748 5906 34804 5908
rect 34748 5854 34750 5906
rect 34750 5854 34802 5906
rect 34802 5854 34804 5906
rect 34748 5852 34804 5854
rect 35980 6748 36036 6804
rect 34972 6412 35028 6468
rect 35532 5852 35588 5908
rect 35084 5794 35140 5796
rect 35084 5742 35086 5794
rect 35086 5742 35138 5794
rect 35138 5742 35140 5794
rect 35084 5740 35140 5742
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35756 5740 35812 5796
rect 35644 5180 35700 5236
rect 34860 5068 34916 5124
rect 35980 5122 36036 5124
rect 35980 5070 35982 5122
rect 35982 5070 36034 5122
rect 36034 5070 36036 5122
rect 35980 5068 36036 5070
rect 35196 5010 35252 5012
rect 35196 4958 35198 5010
rect 35198 4958 35250 5010
rect 35250 4958 35252 5010
rect 35196 4956 35252 4958
rect 35644 4844 35700 4900
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35420 3442 35476 3444
rect 35420 3390 35422 3442
rect 35422 3390 35474 3442
rect 35474 3390 35476 3442
rect 35420 3388 35476 3390
rect 36204 6578 36260 6580
rect 36204 6526 36206 6578
rect 36206 6526 36258 6578
rect 36258 6526 36260 6578
rect 36204 6524 36260 6526
rect 36092 4844 36148 4900
rect 36428 8146 36484 8148
rect 36428 8094 36430 8146
rect 36430 8094 36482 8146
rect 36482 8094 36484 8146
rect 36428 8092 36484 8094
rect 36988 10220 37044 10276
rect 37660 9548 37716 9604
rect 37660 8988 37716 9044
rect 36876 8034 36932 8036
rect 36876 7982 36878 8034
rect 36878 7982 36930 8034
rect 36930 7982 36932 8034
rect 36876 7980 36932 7982
rect 37324 8092 37380 8148
rect 36540 6748 36596 6804
rect 36428 6690 36484 6692
rect 36428 6638 36430 6690
rect 36430 6638 36482 6690
rect 36482 6638 36484 6690
rect 36428 6636 36484 6638
rect 36652 6524 36708 6580
rect 36876 6466 36932 6468
rect 36876 6414 36878 6466
rect 36878 6414 36930 6466
rect 36930 6414 36932 6466
rect 36876 6412 36932 6414
rect 36988 6076 37044 6132
rect 36316 4732 36372 4788
rect 35868 4060 35924 4116
rect 36764 5964 36820 6020
rect 35868 1372 35924 1428
rect 36204 3388 36260 3444
rect 36876 5740 36932 5796
rect 36764 2380 36820 2436
rect 37436 6690 37492 6692
rect 37436 6638 37438 6690
rect 37438 6638 37490 6690
rect 37490 6638 37492 6690
rect 37436 6636 37492 6638
rect 37436 5404 37492 5460
rect 38556 10780 38612 10836
rect 38108 10220 38164 10276
rect 37996 9042 38052 9044
rect 37996 8990 37998 9042
rect 37998 8990 38050 9042
rect 38050 8990 38052 9042
rect 37996 8988 38052 8990
rect 37772 7980 37828 8036
rect 39340 10834 39396 10836
rect 39340 10782 39342 10834
rect 39342 10782 39394 10834
rect 39394 10782 39396 10834
rect 39340 10780 39396 10782
rect 38668 8930 38724 8932
rect 38668 8878 38670 8930
rect 38670 8878 38722 8930
rect 38722 8878 38724 8930
rect 38668 8876 38724 8878
rect 39228 8876 39284 8932
rect 39004 8540 39060 8596
rect 38220 6636 38276 6692
rect 37660 5180 37716 5236
rect 38108 6076 38164 6132
rect 37996 5010 38052 5012
rect 37996 4958 37998 5010
rect 37998 4958 38050 5010
rect 38050 4958 38052 5010
rect 37996 4956 38052 4958
rect 38220 4956 38276 5012
rect 37548 4844 37604 4900
rect 38892 8092 38948 8148
rect 39900 9996 39956 10052
rect 39900 9436 39956 9492
rect 39004 7308 39060 7364
rect 38780 6636 38836 6692
rect 38892 6524 38948 6580
rect 38668 5010 38724 5012
rect 38668 4958 38670 5010
rect 38670 4958 38722 5010
rect 38722 4958 38724 5010
rect 38668 4956 38724 4958
rect 39004 4844 39060 4900
rect 38668 4172 38724 4228
rect 39676 6578 39732 6580
rect 39676 6526 39678 6578
rect 39678 6526 39730 6578
rect 39730 6526 39732 6578
rect 39676 6524 39732 6526
rect 40236 25564 40292 25620
rect 40908 10444 40964 10500
rect 40124 9212 40180 9268
rect 40236 8540 40292 8596
rect 39340 6130 39396 6132
rect 39340 6078 39342 6130
rect 39342 6078 39394 6130
rect 39394 6078 39396 6130
rect 39340 6076 39396 6078
rect 39564 5964 39620 6020
rect 39452 5906 39508 5908
rect 39452 5854 39454 5906
rect 39454 5854 39506 5906
rect 39506 5854 39508 5906
rect 39452 5852 39508 5854
rect 39228 5180 39284 5236
rect 40012 5292 40068 5348
rect 39452 4562 39508 4564
rect 39452 4510 39454 4562
rect 39454 4510 39506 4562
rect 39506 4510 39508 4562
rect 39452 4508 39508 4510
rect 40124 4844 40180 4900
rect 39900 4060 39956 4116
rect 39676 3948 39732 4004
rect 39116 2940 39172 2996
rect 40348 8146 40404 8148
rect 40348 8094 40350 8146
rect 40350 8094 40402 8146
rect 40402 8094 40404 8146
rect 40348 8092 40404 8094
rect 40348 6524 40404 6580
rect 40572 6578 40628 6580
rect 40572 6526 40574 6578
rect 40574 6526 40626 6578
rect 40626 6526 40628 6578
rect 40572 6524 40628 6526
rect 40908 6748 40964 6804
rect 44716 22876 44772 22932
rect 43036 15820 43092 15876
rect 41580 10444 41636 10500
rect 42700 10444 42756 10500
rect 41916 9266 41972 9268
rect 41916 9214 41918 9266
rect 41918 9214 41970 9266
rect 41970 9214 41972 9266
rect 41916 9212 41972 9214
rect 41468 8988 41524 9044
rect 41356 8540 41412 8596
rect 43260 11340 43316 11396
rect 43148 11116 43204 11172
rect 41356 7308 41412 7364
rect 40460 6188 40516 6244
rect 40460 6018 40516 6020
rect 40460 5966 40462 6018
rect 40462 5966 40514 6018
rect 40514 5966 40516 6018
rect 40460 5964 40516 5966
rect 40348 4338 40404 4340
rect 40348 4286 40350 4338
rect 40350 4286 40402 4338
rect 40402 4286 40404 4338
rect 40348 4284 40404 4286
rect 40572 4956 40628 5012
rect 40572 4732 40628 4788
rect 40796 4562 40852 4564
rect 40796 4510 40798 4562
rect 40798 4510 40850 4562
rect 40850 4510 40852 4562
rect 40796 4508 40852 4510
rect 40684 4396 40740 4452
rect 40796 4338 40852 4340
rect 40796 4286 40798 4338
rect 40798 4286 40850 4338
rect 40850 4286 40852 4338
rect 40796 4284 40852 4286
rect 40796 4060 40852 4116
rect 41356 6188 41412 6244
rect 41244 3612 41300 3668
rect 41804 6636 41860 6692
rect 41804 6412 41860 6468
rect 42252 8034 42308 8036
rect 42252 7982 42254 8034
rect 42254 7982 42306 8034
rect 42306 7982 42308 8034
rect 42252 7980 42308 7982
rect 42588 7868 42644 7924
rect 42812 7586 42868 7588
rect 42812 7534 42814 7586
rect 42814 7534 42866 7586
rect 42866 7534 42868 7586
rect 42812 7532 42868 7534
rect 42028 6300 42084 6356
rect 42140 6524 42196 6580
rect 41916 5740 41972 5796
rect 41580 4732 41636 4788
rect 41692 4226 41748 4228
rect 41692 4174 41694 4226
rect 41694 4174 41746 4226
rect 41746 4174 41748 4226
rect 41692 4172 41748 4174
rect 42476 6636 42532 6692
rect 43036 8540 43092 8596
rect 42700 6300 42756 6356
rect 42812 6188 42868 6244
rect 43036 7868 43092 7924
rect 42812 5628 42868 5684
rect 42588 5234 42644 5236
rect 42588 5182 42590 5234
rect 42590 5182 42642 5234
rect 42642 5182 42644 5234
rect 42588 5180 42644 5182
rect 42364 4450 42420 4452
rect 42364 4398 42366 4450
rect 42366 4398 42418 4450
rect 42418 4398 42420 4450
rect 42364 4396 42420 4398
rect 42252 4338 42308 4340
rect 42252 4286 42254 4338
rect 42254 4286 42306 4338
rect 42306 4286 42308 4338
rect 42252 4284 42308 4286
rect 42588 4338 42644 4340
rect 42588 4286 42590 4338
rect 42590 4286 42642 4338
rect 42642 4286 42644 4338
rect 42588 4284 42644 4286
rect 41804 3666 41860 3668
rect 41804 3614 41806 3666
rect 41806 3614 41858 3666
rect 41858 3614 41860 3666
rect 41804 3612 41860 3614
rect 41356 3276 41412 3332
rect 43036 4956 43092 5012
rect 43484 9436 43540 9492
rect 43484 8988 43540 9044
rect 43932 8988 43988 9044
rect 44380 8988 44436 9044
rect 44044 8204 44100 8260
rect 43708 7756 43764 7812
rect 43932 7756 43988 7812
rect 43820 6466 43876 6468
rect 43820 6414 43822 6466
rect 43822 6414 43874 6466
rect 43874 6414 43876 6466
rect 43820 6412 43876 6414
rect 44156 7586 44212 7588
rect 44156 7534 44158 7586
rect 44158 7534 44210 7586
rect 44210 7534 44212 7586
rect 44156 7532 44212 7534
rect 44044 6524 44100 6580
rect 43260 5122 43316 5124
rect 43260 5070 43262 5122
rect 43262 5070 43314 5122
rect 43314 5070 43316 5122
rect 43260 5068 43316 5070
rect 43372 4844 43428 4900
rect 43260 4450 43316 4452
rect 43260 4398 43262 4450
rect 43262 4398 43314 4450
rect 43314 4398 43316 4450
rect 43260 4396 43316 4398
rect 43148 4284 43204 4340
rect 42588 3724 42644 3780
rect 43932 4956 43988 5012
rect 44604 6412 44660 6468
rect 44156 6018 44212 6020
rect 44156 5966 44158 6018
rect 44158 5966 44210 6018
rect 44210 5966 44212 6018
rect 44156 5964 44212 5966
rect 44940 10780 44996 10836
rect 45276 10780 45332 10836
rect 45724 27132 45780 27188
rect 45052 10668 45108 10724
rect 44828 8540 44884 8596
rect 44828 7756 44884 7812
rect 48636 23772 48692 23828
rect 46956 23660 47012 23716
rect 46284 21308 46340 21364
rect 45724 10556 45780 10612
rect 46172 11564 46228 11620
rect 46060 10498 46116 10500
rect 46060 10446 46062 10498
rect 46062 10446 46114 10498
rect 46114 10446 46116 10498
rect 46060 10444 46116 10446
rect 45052 7980 45108 8036
rect 45724 9324 45780 9380
rect 45836 9212 45892 9268
rect 45500 8540 45556 8596
rect 45724 8764 45780 8820
rect 46172 9324 46228 9380
rect 45724 8204 45780 8260
rect 45724 7980 45780 8036
rect 44380 4732 44436 4788
rect 45276 5740 45332 5796
rect 45612 6690 45668 6692
rect 45612 6638 45614 6690
rect 45614 6638 45666 6690
rect 45666 6638 45668 6690
rect 45612 6636 45668 6638
rect 45500 5740 45556 5796
rect 45052 5180 45108 5236
rect 45388 4284 45444 4340
rect 44380 4172 44436 4228
rect 45500 3500 45556 3556
rect 45388 3442 45444 3444
rect 45388 3390 45390 3442
rect 45390 3390 45442 3442
rect 45442 3390 45444 3442
rect 45388 3388 45444 3390
rect 45836 7084 45892 7140
rect 46844 17500 46900 17556
rect 46620 11170 46676 11172
rect 46620 11118 46622 11170
rect 46622 11118 46674 11170
rect 46674 11118 46676 11170
rect 46620 11116 46676 11118
rect 46396 10834 46452 10836
rect 46396 10782 46398 10834
rect 46398 10782 46450 10834
rect 46450 10782 46452 10834
rect 46396 10780 46452 10782
rect 46620 10780 46676 10836
rect 46620 10556 46676 10612
rect 46508 9154 46564 9156
rect 46508 9102 46510 9154
rect 46510 9102 46562 9154
rect 46562 9102 46564 9154
rect 46508 9100 46564 9102
rect 46396 7980 46452 8036
rect 46172 7308 46228 7364
rect 46172 6636 46228 6692
rect 46060 6300 46116 6356
rect 45948 6188 46004 6244
rect 46396 6636 46452 6692
rect 46284 6524 46340 6580
rect 46508 6578 46564 6580
rect 46508 6526 46510 6578
rect 46510 6526 46562 6578
rect 46562 6526 46564 6578
rect 46508 6524 46564 6526
rect 46172 5964 46228 6020
rect 46396 6412 46452 6468
rect 45948 5346 46004 5348
rect 45948 5294 45950 5346
rect 45950 5294 46002 5346
rect 46002 5294 46004 5346
rect 45948 5292 46004 5294
rect 46284 5852 46340 5908
rect 46172 3724 46228 3780
rect 46732 10444 46788 10500
rect 47964 17052 48020 17108
rect 46956 11564 47012 11620
rect 46844 9266 46900 9268
rect 46844 9214 46846 9266
rect 46846 9214 46898 9266
rect 46898 9214 46900 9266
rect 46844 9212 46900 9214
rect 47852 10332 47908 10388
rect 47180 9100 47236 9156
rect 46956 7474 47012 7476
rect 46956 7422 46958 7474
rect 46958 7422 47010 7474
rect 47010 7422 47012 7474
rect 46956 7420 47012 7422
rect 46732 7308 46788 7364
rect 46620 5628 46676 5684
rect 47292 7868 47348 7924
rect 47852 7196 47908 7252
rect 50556 101946 50612 101948
rect 50556 101894 50558 101946
rect 50558 101894 50610 101946
rect 50610 101894 50612 101946
rect 50556 101892 50612 101894
rect 50660 101946 50716 101948
rect 50660 101894 50662 101946
rect 50662 101894 50714 101946
rect 50714 101894 50716 101946
rect 50660 101892 50716 101894
rect 50764 101946 50820 101948
rect 50764 101894 50766 101946
rect 50766 101894 50818 101946
rect 50818 101894 50820 101946
rect 50764 101892 50820 101894
rect 50556 100378 50612 100380
rect 50556 100326 50558 100378
rect 50558 100326 50610 100378
rect 50610 100326 50612 100378
rect 50556 100324 50612 100326
rect 50660 100378 50716 100380
rect 50660 100326 50662 100378
rect 50662 100326 50714 100378
rect 50714 100326 50716 100378
rect 50660 100324 50716 100326
rect 50764 100378 50820 100380
rect 50764 100326 50766 100378
rect 50766 100326 50818 100378
rect 50818 100326 50820 100378
rect 50764 100324 50820 100326
rect 50556 98810 50612 98812
rect 50556 98758 50558 98810
rect 50558 98758 50610 98810
rect 50610 98758 50612 98810
rect 50556 98756 50612 98758
rect 50660 98810 50716 98812
rect 50660 98758 50662 98810
rect 50662 98758 50714 98810
rect 50714 98758 50716 98810
rect 50660 98756 50716 98758
rect 50764 98810 50820 98812
rect 50764 98758 50766 98810
rect 50766 98758 50818 98810
rect 50818 98758 50820 98810
rect 50764 98756 50820 98758
rect 50556 97242 50612 97244
rect 50556 97190 50558 97242
rect 50558 97190 50610 97242
rect 50610 97190 50612 97242
rect 50556 97188 50612 97190
rect 50660 97242 50716 97244
rect 50660 97190 50662 97242
rect 50662 97190 50714 97242
rect 50714 97190 50716 97242
rect 50660 97188 50716 97190
rect 50764 97242 50820 97244
rect 50764 97190 50766 97242
rect 50766 97190 50818 97242
rect 50818 97190 50820 97242
rect 50764 97188 50820 97190
rect 50556 95674 50612 95676
rect 50556 95622 50558 95674
rect 50558 95622 50610 95674
rect 50610 95622 50612 95674
rect 50556 95620 50612 95622
rect 50660 95674 50716 95676
rect 50660 95622 50662 95674
rect 50662 95622 50714 95674
rect 50714 95622 50716 95674
rect 50660 95620 50716 95622
rect 50764 95674 50820 95676
rect 50764 95622 50766 95674
rect 50766 95622 50818 95674
rect 50818 95622 50820 95674
rect 50764 95620 50820 95622
rect 50556 94106 50612 94108
rect 50556 94054 50558 94106
rect 50558 94054 50610 94106
rect 50610 94054 50612 94106
rect 50556 94052 50612 94054
rect 50660 94106 50716 94108
rect 50660 94054 50662 94106
rect 50662 94054 50714 94106
rect 50714 94054 50716 94106
rect 50660 94052 50716 94054
rect 50764 94106 50820 94108
rect 50764 94054 50766 94106
rect 50766 94054 50818 94106
rect 50818 94054 50820 94106
rect 50764 94052 50820 94054
rect 50556 92538 50612 92540
rect 50556 92486 50558 92538
rect 50558 92486 50610 92538
rect 50610 92486 50612 92538
rect 50556 92484 50612 92486
rect 50660 92538 50716 92540
rect 50660 92486 50662 92538
rect 50662 92486 50714 92538
rect 50714 92486 50716 92538
rect 50660 92484 50716 92486
rect 50764 92538 50820 92540
rect 50764 92486 50766 92538
rect 50766 92486 50818 92538
rect 50818 92486 50820 92538
rect 50764 92484 50820 92486
rect 50556 90970 50612 90972
rect 50556 90918 50558 90970
rect 50558 90918 50610 90970
rect 50610 90918 50612 90970
rect 50556 90916 50612 90918
rect 50660 90970 50716 90972
rect 50660 90918 50662 90970
rect 50662 90918 50714 90970
rect 50714 90918 50716 90970
rect 50660 90916 50716 90918
rect 50764 90970 50820 90972
rect 50764 90918 50766 90970
rect 50766 90918 50818 90970
rect 50818 90918 50820 90970
rect 50764 90916 50820 90918
rect 50556 89402 50612 89404
rect 50556 89350 50558 89402
rect 50558 89350 50610 89402
rect 50610 89350 50612 89402
rect 50556 89348 50612 89350
rect 50660 89402 50716 89404
rect 50660 89350 50662 89402
rect 50662 89350 50714 89402
rect 50714 89350 50716 89402
rect 50660 89348 50716 89350
rect 50764 89402 50820 89404
rect 50764 89350 50766 89402
rect 50766 89350 50818 89402
rect 50818 89350 50820 89402
rect 50764 89348 50820 89350
rect 50556 87834 50612 87836
rect 50556 87782 50558 87834
rect 50558 87782 50610 87834
rect 50610 87782 50612 87834
rect 50556 87780 50612 87782
rect 50660 87834 50716 87836
rect 50660 87782 50662 87834
rect 50662 87782 50714 87834
rect 50714 87782 50716 87834
rect 50660 87780 50716 87782
rect 50764 87834 50820 87836
rect 50764 87782 50766 87834
rect 50766 87782 50818 87834
rect 50818 87782 50820 87834
rect 50764 87780 50820 87782
rect 50556 86266 50612 86268
rect 50556 86214 50558 86266
rect 50558 86214 50610 86266
rect 50610 86214 50612 86266
rect 50556 86212 50612 86214
rect 50660 86266 50716 86268
rect 50660 86214 50662 86266
rect 50662 86214 50714 86266
rect 50714 86214 50716 86266
rect 50660 86212 50716 86214
rect 50764 86266 50820 86268
rect 50764 86214 50766 86266
rect 50766 86214 50818 86266
rect 50818 86214 50820 86266
rect 50764 86212 50820 86214
rect 50556 84698 50612 84700
rect 50556 84646 50558 84698
rect 50558 84646 50610 84698
rect 50610 84646 50612 84698
rect 50556 84644 50612 84646
rect 50660 84698 50716 84700
rect 50660 84646 50662 84698
rect 50662 84646 50714 84698
rect 50714 84646 50716 84698
rect 50660 84644 50716 84646
rect 50764 84698 50820 84700
rect 50764 84646 50766 84698
rect 50766 84646 50818 84698
rect 50818 84646 50820 84698
rect 50764 84644 50820 84646
rect 50556 83130 50612 83132
rect 50556 83078 50558 83130
rect 50558 83078 50610 83130
rect 50610 83078 50612 83130
rect 50556 83076 50612 83078
rect 50660 83130 50716 83132
rect 50660 83078 50662 83130
rect 50662 83078 50714 83130
rect 50714 83078 50716 83130
rect 50660 83076 50716 83078
rect 50764 83130 50820 83132
rect 50764 83078 50766 83130
rect 50766 83078 50818 83130
rect 50818 83078 50820 83130
rect 50764 83076 50820 83078
rect 50556 81562 50612 81564
rect 50556 81510 50558 81562
rect 50558 81510 50610 81562
rect 50610 81510 50612 81562
rect 50556 81508 50612 81510
rect 50660 81562 50716 81564
rect 50660 81510 50662 81562
rect 50662 81510 50714 81562
rect 50714 81510 50716 81562
rect 50660 81508 50716 81510
rect 50764 81562 50820 81564
rect 50764 81510 50766 81562
rect 50766 81510 50818 81562
rect 50818 81510 50820 81562
rect 50764 81508 50820 81510
rect 50556 79994 50612 79996
rect 50556 79942 50558 79994
rect 50558 79942 50610 79994
rect 50610 79942 50612 79994
rect 50556 79940 50612 79942
rect 50660 79994 50716 79996
rect 50660 79942 50662 79994
rect 50662 79942 50714 79994
rect 50714 79942 50716 79994
rect 50660 79940 50716 79942
rect 50764 79994 50820 79996
rect 50764 79942 50766 79994
rect 50766 79942 50818 79994
rect 50818 79942 50820 79994
rect 50764 79940 50820 79942
rect 50556 78426 50612 78428
rect 50556 78374 50558 78426
rect 50558 78374 50610 78426
rect 50610 78374 50612 78426
rect 50556 78372 50612 78374
rect 50660 78426 50716 78428
rect 50660 78374 50662 78426
rect 50662 78374 50714 78426
rect 50714 78374 50716 78426
rect 50660 78372 50716 78374
rect 50764 78426 50820 78428
rect 50764 78374 50766 78426
rect 50766 78374 50818 78426
rect 50818 78374 50820 78426
rect 50764 78372 50820 78374
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 48748 20972 48804 21028
rect 49196 30268 49252 30324
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 52780 25452 52836 25508
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 48972 16940 49028 16996
rect 48636 10332 48692 10388
rect 48300 9100 48356 9156
rect 47628 6748 47684 6804
rect 47740 6636 47796 6692
rect 47628 6188 47684 6244
rect 47628 6018 47684 6020
rect 47628 5966 47630 6018
rect 47630 5966 47682 6018
rect 47682 5966 47684 6018
rect 47628 5964 47684 5966
rect 47404 5906 47460 5908
rect 47404 5854 47406 5906
rect 47406 5854 47458 5906
rect 47458 5854 47460 5906
rect 47404 5852 47460 5854
rect 46844 3554 46900 3556
rect 46844 3502 46846 3554
rect 46846 3502 46898 3554
rect 46898 3502 46900 3554
rect 46844 3500 46900 3502
rect 46284 3276 46340 3332
rect 48188 6412 48244 6468
rect 48076 6076 48132 6132
rect 47964 5740 48020 5796
rect 47852 5628 47908 5684
rect 48636 9154 48692 9156
rect 48636 9102 48638 9154
rect 48638 9102 48690 9154
rect 48690 9102 48692 9154
rect 48636 9100 48692 9102
rect 48972 9212 49028 9268
rect 49084 9996 49140 10052
rect 48412 7362 48468 7364
rect 48412 7310 48414 7362
rect 48414 7310 48466 7362
rect 48466 7310 48468 7362
rect 48412 7308 48468 7310
rect 48636 7196 48692 7252
rect 48748 7420 48804 7476
rect 48412 4338 48468 4340
rect 48412 4286 48414 4338
rect 48414 4286 48466 4338
rect 48466 4286 48468 4338
rect 48412 4284 48468 4286
rect 47740 3442 47796 3444
rect 47740 3390 47742 3442
rect 47742 3390 47794 3442
rect 47794 3390 47796 3442
rect 47740 3388 47796 3390
rect 48972 6578 49028 6580
rect 48972 6526 48974 6578
rect 48974 6526 49026 6578
rect 49026 6526 49028 6578
rect 48972 6524 49028 6526
rect 48972 6300 49028 6356
rect 48860 6018 48916 6020
rect 48860 5966 48862 6018
rect 48862 5966 48914 6018
rect 48914 5966 48916 6018
rect 48860 5964 48916 5966
rect 49084 5404 49140 5460
rect 48860 5010 48916 5012
rect 48860 4958 48862 5010
rect 48862 4958 48914 5010
rect 48914 4958 48916 5010
rect 48860 4956 48916 4958
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 51548 12460 51604 12516
rect 51100 11282 51156 11284
rect 51100 11230 51102 11282
rect 51102 11230 51154 11282
rect 51154 11230 51156 11282
rect 51100 11228 51156 11230
rect 51324 11228 51380 11284
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 51100 10780 51156 10836
rect 50876 10556 50932 10612
rect 49868 10498 49924 10500
rect 49868 10446 49870 10498
rect 49870 10446 49922 10498
rect 49922 10446 49924 10498
rect 49868 10444 49924 10446
rect 49532 9100 49588 9156
rect 49980 8988 50036 9044
rect 49756 7308 49812 7364
rect 49644 6412 49700 6468
rect 50316 9042 50372 9044
rect 50316 8990 50318 9042
rect 50318 8990 50370 9042
rect 50370 8990 50372 9042
rect 50316 8988 50372 8990
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50428 6972 50484 7028
rect 50988 7868 51044 7924
rect 51212 9996 51268 10052
rect 51996 11788 52052 11844
rect 51660 11170 51716 11172
rect 51660 11118 51662 11170
rect 51662 11118 51714 11170
rect 51714 11118 51716 11170
rect 51660 11116 51716 11118
rect 51884 10556 51940 10612
rect 51212 6972 51268 7028
rect 50876 6636 50932 6692
rect 51548 9660 51604 9716
rect 52892 23548 52948 23604
rect 53564 23548 53620 23604
rect 58156 21420 58212 21476
rect 57036 19068 57092 19124
rect 55804 14588 55860 14644
rect 52892 11788 52948 11844
rect 52780 11170 52836 11172
rect 52780 11118 52782 11170
rect 52782 11118 52834 11170
rect 52834 11118 52836 11170
rect 52780 11116 52836 11118
rect 51324 6524 51380 6580
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 49980 5964 50036 6020
rect 51212 5292 51268 5348
rect 49756 5234 49812 5236
rect 49756 5182 49758 5234
rect 49758 5182 49810 5234
rect 49810 5182 49812 5234
rect 49756 5180 49812 5182
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50876 4172 50932 4228
rect 49644 3388 49700 3444
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 51436 5180 51492 5236
rect 51884 7980 51940 8036
rect 52668 10556 52724 10612
rect 52332 9996 52388 10052
rect 52444 8764 52500 8820
rect 53564 10444 53620 10500
rect 53676 9938 53732 9940
rect 53676 9886 53678 9938
rect 53678 9886 53730 9938
rect 53730 9886 53732 9938
rect 53676 9884 53732 9886
rect 52780 8764 52836 8820
rect 53340 8764 53396 8820
rect 52556 8204 52612 8260
rect 54684 10332 54740 10388
rect 52332 8034 52388 8036
rect 52332 7982 52334 8034
rect 52334 7982 52386 8034
rect 52386 7982 52388 8034
rect 52332 7980 52388 7982
rect 52220 7868 52276 7924
rect 52108 6748 52164 6804
rect 51996 4620 52052 4676
rect 51996 4284 52052 4340
rect 52220 6636 52276 6692
rect 53452 6690 53508 6692
rect 53452 6638 53454 6690
rect 53454 6638 53506 6690
rect 53506 6638 53508 6690
rect 53452 6636 53508 6638
rect 52332 6578 52388 6580
rect 52332 6526 52334 6578
rect 52334 6526 52386 6578
rect 52386 6526 52388 6578
rect 52332 6524 52388 6526
rect 52108 2828 52164 2884
rect 52444 5628 52500 5684
rect 53788 6748 53844 6804
rect 53900 9884 53956 9940
rect 55468 11116 55524 11172
rect 55020 9884 55076 9940
rect 55020 9212 55076 9268
rect 53900 8988 53956 9044
rect 54796 8988 54852 9044
rect 54012 8258 54068 8260
rect 54012 8206 54014 8258
rect 54014 8206 54066 8258
rect 54066 8206 54068 8258
rect 54012 8204 54068 8206
rect 53564 5292 53620 5348
rect 52556 5122 52612 5124
rect 52556 5070 52558 5122
rect 52558 5070 52610 5122
rect 52610 5070 52612 5122
rect 52556 5068 52612 5070
rect 53788 5122 53844 5124
rect 53788 5070 53790 5122
rect 53790 5070 53842 5122
rect 53842 5070 53844 5122
rect 53788 5068 53844 5070
rect 54236 7980 54292 8036
rect 54796 6188 54852 6244
rect 55244 9100 55300 9156
rect 55468 9100 55524 9156
rect 55356 7474 55412 7476
rect 55356 7422 55358 7474
rect 55358 7422 55410 7474
rect 55410 7422 55412 7474
rect 55356 7420 55412 7422
rect 55244 6412 55300 6468
rect 54012 4956 54068 5012
rect 55692 9548 55748 9604
rect 55692 8988 55748 9044
rect 56588 13916 56644 13972
rect 56252 12460 56308 12516
rect 56140 11564 56196 11620
rect 56028 11170 56084 11172
rect 56028 11118 56030 11170
rect 56030 11118 56082 11170
rect 56082 11118 56084 11170
rect 56028 11116 56084 11118
rect 55916 10556 55972 10612
rect 56028 10332 56084 10388
rect 56140 10444 56196 10500
rect 56140 9042 56196 9044
rect 56140 8990 56142 9042
rect 56142 8990 56194 9042
rect 56194 8990 56196 9042
rect 56140 8988 56196 8990
rect 56476 10498 56532 10500
rect 56476 10446 56478 10498
rect 56478 10446 56530 10498
rect 56530 10446 56532 10498
rect 56476 10444 56532 10446
rect 56364 9548 56420 9604
rect 55916 8034 55972 8036
rect 55916 7982 55918 8034
rect 55918 7982 55970 8034
rect 55970 7982 55972 8034
rect 55916 7980 55972 7982
rect 55580 7420 55636 7476
rect 55804 7420 55860 7476
rect 55692 6018 55748 6020
rect 55692 5966 55694 6018
rect 55694 5966 55746 6018
rect 55746 5966 55748 6018
rect 55692 5964 55748 5966
rect 54572 5234 54628 5236
rect 54572 5182 54574 5234
rect 54574 5182 54626 5234
rect 54626 5182 54628 5234
rect 54572 5180 54628 5182
rect 54684 4172 54740 4228
rect 55580 4226 55636 4228
rect 55580 4174 55582 4226
rect 55582 4174 55634 4226
rect 55634 4174 55636 4226
rect 55580 4172 55636 4174
rect 55020 3442 55076 3444
rect 55020 3390 55022 3442
rect 55022 3390 55074 3442
rect 55074 3390 55076 3442
rect 55020 3388 55076 3390
rect 57036 12460 57092 12516
rect 57708 15932 57764 15988
rect 57372 12290 57428 12292
rect 57372 12238 57374 12290
rect 57374 12238 57426 12290
rect 57426 12238 57428 12290
rect 57372 12236 57428 12238
rect 56812 10556 56868 10612
rect 56924 10668 56980 10724
rect 56700 9042 56756 9044
rect 56700 8990 56702 9042
rect 56702 8990 56754 9042
rect 56754 8990 56756 9042
rect 56700 8988 56756 8990
rect 57036 7644 57092 7700
rect 56588 6524 56644 6580
rect 56364 5964 56420 6020
rect 56700 5964 56756 6020
rect 57148 7084 57204 7140
rect 57148 6690 57204 6692
rect 57148 6638 57150 6690
rect 57150 6638 57202 6690
rect 57202 6638 57204 6690
rect 57148 6636 57204 6638
rect 57036 5068 57092 5124
rect 57484 10722 57540 10724
rect 57484 10670 57486 10722
rect 57486 10670 57538 10722
rect 57538 10670 57540 10722
rect 57484 10668 57540 10670
rect 57484 7644 57540 7700
rect 57932 12460 57988 12516
rect 57484 6018 57540 6020
rect 57484 5966 57486 6018
rect 57486 5966 57538 6018
rect 57538 5966 57540 6018
rect 57484 5964 57540 5966
rect 57148 4956 57204 5012
rect 56364 3388 56420 3444
rect 57484 4338 57540 4340
rect 57484 4286 57486 4338
rect 57486 4286 57538 4338
rect 57538 4286 57540 4338
rect 57484 4284 57540 4286
rect 57708 6018 57764 6020
rect 57708 5966 57710 6018
rect 57710 5966 57762 6018
rect 57762 5966 57764 6018
rect 57708 5964 57764 5966
rect 57932 7084 57988 7140
rect 58044 6578 58100 6580
rect 58044 6526 58046 6578
rect 58046 6526 58098 6578
rect 58098 6526 58100 6578
rect 58044 6524 58100 6526
rect 57932 5180 57988 5236
rect 57708 4620 57764 4676
rect 65916 116842 65972 116844
rect 65916 116790 65918 116842
rect 65918 116790 65970 116842
rect 65970 116790 65972 116842
rect 65916 116788 65972 116790
rect 66020 116842 66076 116844
rect 66020 116790 66022 116842
rect 66022 116790 66074 116842
rect 66074 116790 66076 116842
rect 66020 116788 66076 116790
rect 66124 116842 66180 116844
rect 66124 116790 66126 116842
rect 66126 116790 66178 116842
rect 66178 116790 66180 116842
rect 66124 116788 66180 116790
rect 73052 116508 73108 116564
rect 67116 116172 67172 116228
rect 67564 116226 67620 116228
rect 67564 116174 67566 116226
rect 67566 116174 67618 116226
rect 67618 116174 67620 116226
rect 67564 116172 67620 116174
rect 63196 115554 63252 115556
rect 63196 115502 63198 115554
rect 63198 115502 63250 115554
rect 63250 115502 63252 115554
rect 63196 115500 63252 115502
rect 63756 115500 63812 115556
rect 69916 116172 69972 116228
rect 67900 115554 67956 115556
rect 67900 115502 67902 115554
rect 67902 115502 67954 115554
rect 67954 115502 67956 115554
rect 67900 115500 67956 115502
rect 68572 115500 68628 115556
rect 65916 115274 65972 115276
rect 65916 115222 65918 115274
rect 65918 115222 65970 115274
rect 65970 115222 65972 115274
rect 65916 115220 65972 115222
rect 66020 115274 66076 115276
rect 66020 115222 66022 115274
rect 66022 115222 66074 115274
rect 66074 115222 66076 115274
rect 66020 115220 66076 115222
rect 66124 115274 66180 115276
rect 66124 115222 66126 115274
rect 66126 115222 66178 115274
rect 66178 115222 66180 115274
rect 66124 115220 66180 115222
rect 64204 115052 64260 115108
rect 64988 115052 65044 115108
rect 65916 113706 65972 113708
rect 65916 113654 65918 113706
rect 65918 113654 65970 113706
rect 65970 113654 65972 113706
rect 65916 113652 65972 113654
rect 66020 113706 66076 113708
rect 66020 113654 66022 113706
rect 66022 113654 66074 113706
rect 66074 113654 66076 113706
rect 66020 113652 66076 113654
rect 66124 113706 66180 113708
rect 66124 113654 66126 113706
rect 66126 113654 66178 113706
rect 66178 113654 66180 113706
rect 66124 113652 66180 113654
rect 65916 112138 65972 112140
rect 65916 112086 65918 112138
rect 65918 112086 65970 112138
rect 65970 112086 65972 112138
rect 65916 112084 65972 112086
rect 66020 112138 66076 112140
rect 66020 112086 66022 112138
rect 66022 112086 66074 112138
rect 66074 112086 66076 112138
rect 66020 112084 66076 112086
rect 66124 112138 66180 112140
rect 66124 112086 66126 112138
rect 66126 112086 66178 112138
rect 66178 112086 66180 112138
rect 66124 112084 66180 112086
rect 65916 110570 65972 110572
rect 65916 110518 65918 110570
rect 65918 110518 65970 110570
rect 65970 110518 65972 110570
rect 65916 110516 65972 110518
rect 66020 110570 66076 110572
rect 66020 110518 66022 110570
rect 66022 110518 66074 110570
rect 66074 110518 66076 110570
rect 66020 110516 66076 110518
rect 66124 110570 66180 110572
rect 66124 110518 66126 110570
rect 66126 110518 66178 110570
rect 66178 110518 66180 110570
rect 66124 110516 66180 110518
rect 65916 109002 65972 109004
rect 65916 108950 65918 109002
rect 65918 108950 65970 109002
rect 65970 108950 65972 109002
rect 65916 108948 65972 108950
rect 66020 109002 66076 109004
rect 66020 108950 66022 109002
rect 66022 108950 66074 109002
rect 66074 108950 66076 109002
rect 66020 108948 66076 108950
rect 66124 109002 66180 109004
rect 66124 108950 66126 109002
rect 66126 108950 66178 109002
rect 66178 108950 66180 109002
rect 66124 108948 66180 108950
rect 65916 107434 65972 107436
rect 65916 107382 65918 107434
rect 65918 107382 65970 107434
rect 65970 107382 65972 107434
rect 65916 107380 65972 107382
rect 66020 107434 66076 107436
rect 66020 107382 66022 107434
rect 66022 107382 66074 107434
rect 66074 107382 66076 107434
rect 66020 107380 66076 107382
rect 66124 107434 66180 107436
rect 66124 107382 66126 107434
rect 66126 107382 66178 107434
rect 66178 107382 66180 107434
rect 66124 107380 66180 107382
rect 65916 105866 65972 105868
rect 65916 105814 65918 105866
rect 65918 105814 65970 105866
rect 65970 105814 65972 105866
rect 65916 105812 65972 105814
rect 66020 105866 66076 105868
rect 66020 105814 66022 105866
rect 66022 105814 66074 105866
rect 66074 105814 66076 105866
rect 66020 105812 66076 105814
rect 66124 105866 66180 105868
rect 66124 105814 66126 105866
rect 66126 105814 66178 105866
rect 66178 105814 66180 105866
rect 66124 105812 66180 105814
rect 65916 104298 65972 104300
rect 65916 104246 65918 104298
rect 65918 104246 65970 104298
rect 65970 104246 65972 104298
rect 65916 104244 65972 104246
rect 66020 104298 66076 104300
rect 66020 104246 66022 104298
rect 66022 104246 66074 104298
rect 66074 104246 66076 104298
rect 66020 104244 66076 104246
rect 66124 104298 66180 104300
rect 66124 104246 66126 104298
rect 66126 104246 66178 104298
rect 66178 104246 66180 104298
rect 66124 104244 66180 104246
rect 65916 102730 65972 102732
rect 65916 102678 65918 102730
rect 65918 102678 65970 102730
rect 65970 102678 65972 102730
rect 65916 102676 65972 102678
rect 66020 102730 66076 102732
rect 66020 102678 66022 102730
rect 66022 102678 66074 102730
rect 66074 102678 66076 102730
rect 66020 102676 66076 102678
rect 66124 102730 66180 102732
rect 66124 102678 66126 102730
rect 66126 102678 66178 102730
rect 66178 102678 66180 102730
rect 66124 102676 66180 102678
rect 65916 101162 65972 101164
rect 65916 101110 65918 101162
rect 65918 101110 65970 101162
rect 65970 101110 65972 101162
rect 65916 101108 65972 101110
rect 66020 101162 66076 101164
rect 66020 101110 66022 101162
rect 66022 101110 66074 101162
rect 66074 101110 66076 101162
rect 66020 101108 66076 101110
rect 66124 101162 66180 101164
rect 66124 101110 66126 101162
rect 66126 101110 66178 101162
rect 66178 101110 66180 101162
rect 66124 101108 66180 101110
rect 65916 99594 65972 99596
rect 65916 99542 65918 99594
rect 65918 99542 65970 99594
rect 65970 99542 65972 99594
rect 65916 99540 65972 99542
rect 66020 99594 66076 99596
rect 66020 99542 66022 99594
rect 66022 99542 66074 99594
rect 66074 99542 66076 99594
rect 66020 99540 66076 99542
rect 66124 99594 66180 99596
rect 66124 99542 66126 99594
rect 66126 99542 66178 99594
rect 66178 99542 66180 99594
rect 66124 99540 66180 99542
rect 65916 98026 65972 98028
rect 65916 97974 65918 98026
rect 65918 97974 65970 98026
rect 65970 97974 65972 98026
rect 65916 97972 65972 97974
rect 66020 98026 66076 98028
rect 66020 97974 66022 98026
rect 66022 97974 66074 98026
rect 66074 97974 66076 98026
rect 66020 97972 66076 97974
rect 66124 98026 66180 98028
rect 66124 97974 66126 98026
rect 66126 97974 66178 98026
rect 66178 97974 66180 98026
rect 66124 97972 66180 97974
rect 65916 96458 65972 96460
rect 65916 96406 65918 96458
rect 65918 96406 65970 96458
rect 65970 96406 65972 96458
rect 65916 96404 65972 96406
rect 66020 96458 66076 96460
rect 66020 96406 66022 96458
rect 66022 96406 66074 96458
rect 66074 96406 66076 96458
rect 66020 96404 66076 96406
rect 66124 96458 66180 96460
rect 66124 96406 66126 96458
rect 66126 96406 66178 96458
rect 66178 96406 66180 96458
rect 66124 96404 66180 96406
rect 65916 94890 65972 94892
rect 65916 94838 65918 94890
rect 65918 94838 65970 94890
rect 65970 94838 65972 94890
rect 65916 94836 65972 94838
rect 66020 94890 66076 94892
rect 66020 94838 66022 94890
rect 66022 94838 66074 94890
rect 66074 94838 66076 94890
rect 66020 94836 66076 94838
rect 66124 94890 66180 94892
rect 66124 94838 66126 94890
rect 66126 94838 66178 94890
rect 66178 94838 66180 94890
rect 66124 94836 66180 94838
rect 65916 93322 65972 93324
rect 65916 93270 65918 93322
rect 65918 93270 65970 93322
rect 65970 93270 65972 93322
rect 65916 93268 65972 93270
rect 66020 93322 66076 93324
rect 66020 93270 66022 93322
rect 66022 93270 66074 93322
rect 66074 93270 66076 93322
rect 66020 93268 66076 93270
rect 66124 93322 66180 93324
rect 66124 93270 66126 93322
rect 66126 93270 66178 93322
rect 66178 93270 66180 93322
rect 66124 93268 66180 93270
rect 65916 91754 65972 91756
rect 65916 91702 65918 91754
rect 65918 91702 65970 91754
rect 65970 91702 65972 91754
rect 65916 91700 65972 91702
rect 66020 91754 66076 91756
rect 66020 91702 66022 91754
rect 66022 91702 66074 91754
rect 66074 91702 66076 91754
rect 66020 91700 66076 91702
rect 66124 91754 66180 91756
rect 66124 91702 66126 91754
rect 66126 91702 66178 91754
rect 66178 91702 66180 91754
rect 66124 91700 66180 91702
rect 65916 90186 65972 90188
rect 65916 90134 65918 90186
rect 65918 90134 65970 90186
rect 65970 90134 65972 90186
rect 65916 90132 65972 90134
rect 66020 90186 66076 90188
rect 66020 90134 66022 90186
rect 66022 90134 66074 90186
rect 66074 90134 66076 90186
rect 66020 90132 66076 90134
rect 66124 90186 66180 90188
rect 66124 90134 66126 90186
rect 66126 90134 66178 90186
rect 66178 90134 66180 90186
rect 66124 90132 66180 90134
rect 65916 88618 65972 88620
rect 65916 88566 65918 88618
rect 65918 88566 65970 88618
rect 65970 88566 65972 88618
rect 65916 88564 65972 88566
rect 66020 88618 66076 88620
rect 66020 88566 66022 88618
rect 66022 88566 66074 88618
rect 66074 88566 66076 88618
rect 66020 88564 66076 88566
rect 66124 88618 66180 88620
rect 66124 88566 66126 88618
rect 66126 88566 66178 88618
rect 66178 88566 66180 88618
rect 66124 88564 66180 88566
rect 65916 87050 65972 87052
rect 65916 86998 65918 87050
rect 65918 86998 65970 87050
rect 65970 86998 65972 87050
rect 65916 86996 65972 86998
rect 66020 87050 66076 87052
rect 66020 86998 66022 87050
rect 66022 86998 66074 87050
rect 66074 86998 66076 87050
rect 66020 86996 66076 86998
rect 66124 87050 66180 87052
rect 66124 86998 66126 87050
rect 66126 86998 66178 87050
rect 66178 86998 66180 87050
rect 66124 86996 66180 86998
rect 65916 85482 65972 85484
rect 65916 85430 65918 85482
rect 65918 85430 65970 85482
rect 65970 85430 65972 85482
rect 65916 85428 65972 85430
rect 66020 85482 66076 85484
rect 66020 85430 66022 85482
rect 66022 85430 66074 85482
rect 66074 85430 66076 85482
rect 66020 85428 66076 85430
rect 66124 85482 66180 85484
rect 66124 85430 66126 85482
rect 66126 85430 66178 85482
rect 66178 85430 66180 85482
rect 66124 85428 66180 85430
rect 65916 83914 65972 83916
rect 65916 83862 65918 83914
rect 65918 83862 65970 83914
rect 65970 83862 65972 83914
rect 65916 83860 65972 83862
rect 66020 83914 66076 83916
rect 66020 83862 66022 83914
rect 66022 83862 66074 83914
rect 66074 83862 66076 83914
rect 66020 83860 66076 83862
rect 66124 83914 66180 83916
rect 66124 83862 66126 83914
rect 66126 83862 66178 83914
rect 66178 83862 66180 83914
rect 66124 83860 66180 83862
rect 65916 82346 65972 82348
rect 65916 82294 65918 82346
rect 65918 82294 65970 82346
rect 65970 82294 65972 82346
rect 65916 82292 65972 82294
rect 66020 82346 66076 82348
rect 66020 82294 66022 82346
rect 66022 82294 66074 82346
rect 66074 82294 66076 82346
rect 66020 82292 66076 82294
rect 66124 82346 66180 82348
rect 66124 82294 66126 82346
rect 66126 82294 66178 82346
rect 66178 82294 66180 82346
rect 66124 82292 66180 82294
rect 65916 80778 65972 80780
rect 65916 80726 65918 80778
rect 65918 80726 65970 80778
rect 65970 80726 65972 80778
rect 65916 80724 65972 80726
rect 66020 80778 66076 80780
rect 66020 80726 66022 80778
rect 66022 80726 66074 80778
rect 66074 80726 66076 80778
rect 66020 80724 66076 80726
rect 66124 80778 66180 80780
rect 66124 80726 66126 80778
rect 66126 80726 66178 80778
rect 66178 80726 66180 80778
rect 66124 80724 66180 80726
rect 65916 79210 65972 79212
rect 65916 79158 65918 79210
rect 65918 79158 65970 79210
rect 65970 79158 65972 79210
rect 65916 79156 65972 79158
rect 66020 79210 66076 79212
rect 66020 79158 66022 79210
rect 66022 79158 66074 79210
rect 66074 79158 66076 79210
rect 66020 79156 66076 79158
rect 66124 79210 66180 79212
rect 66124 79158 66126 79210
rect 66126 79158 66178 79210
rect 66178 79158 66180 79210
rect 66124 79156 66180 79158
rect 65916 77642 65972 77644
rect 65916 77590 65918 77642
rect 65918 77590 65970 77642
rect 65970 77590 65972 77642
rect 65916 77588 65972 77590
rect 66020 77642 66076 77644
rect 66020 77590 66022 77642
rect 66022 77590 66074 77642
rect 66074 77590 66076 77642
rect 66020 77588 66076 77590
rect 66124 77642 66180 77644
rect 66124 77590 66126 77642
rect 66126 77590 66178 77642
rect 66178 77590 66180 77642
rect 66124 77588 66180 77590
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 67900 27356 67956 27412
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 62860 19404 62916 19460
rect 65548 24108 65604 24164
rect 63756 19292 63812 19348
rect 58492 18956 58548 19012
rect 62188 17388 62244 17444
rect 58940 16156 58996 16212
rect 58604 12236 58660 12292
rect 58268 8930 58324 8932
rect 58268 8878 58270 8930
rect 58270 8878 58322 8930
rect 58322 8878 58324 8930
rect 58268 8876 58324 8878
rect 58492 9100 58548 9156
rect 58380 8034 58436 8036
rect 58380 7982 58382 8034
rect 58382 7982 58434 8034
rect 58434 7982 58436 8034
rect 58380 7980 58436 7982
rect 58604 8988 58660 9044
rect 58828 9154 58884 9156
rect 58828 9102 58830 9154
rect 58830 9102 58882 9154
rect 58882 9102 58884 9154
rect 58828 9100 58884 9102
rect 58716 7980 58772 8036
rect 61740 14700 61796 14756
rect 60508 14476 60564 14532
rect 59612 12290 59668 12292
rect 59612 12238 59614 12290
rect 59614 12238 59666 12290
rect 59666 12238 59668 12290
rect 59612 12236 59668 12238
rect 59164 12066 59220 12068
rect 59164 12014 59166 12066
rect 59166 12014 59218 12066
rect 59218 12014 59220 12066
rect 59164 12012 59220 12014
rect 59388 11452 59444 11508
rect 59052 9100 59108 9156
rect 59276 8428 59332 8484
rect 59948 11506 60004 11508
rect 59948 11454 59950 11506
rect 59950 11454 60002 11506
rect 60002 11454 60004 11506
rect 59948 11452 60004 11454
rect 61516 13580 61572 13636
rect 60844 12290 60900 12292
rect 60844 12238 60846 12290
rect 60846 12238 60898 12290
rect 60898 12238 60900 12290
rect 60844 12236 60900 12238
rect 61180 12012 61236 12068
rect 60620 11954 60676 11956
rect 60620 11902 60622 11954
rect 60622 11902 60674 11954
rect 60674 11902 60676 11954
rect 60620 11900 60676 11902
rect 60508 11452 60564 11508
rect 60508 10556 60564 10612
rect 59612 9154 59668 9156
rect 59612 9102 59614 9154
rect 59614 9102 59666 9154
rect 59666 9102 59668 9154
rect 59612 9100 59668 9102
rect 60620 9042 60676 9044
rect 60620 8990 60622 9042
rect 60622 8990 60674 9042
rect 60674 8990 60676 9042
rect 60620 8988 60676 8990
rect 59276 8258 59332 8260
rect 59276 8206 59278 8258
rect 59278 8206 59330 8258
rect 59330 8206 59332 8258
rect 59276 8204 59332 8206
rect 58940 8034 58996 8036
rect 58940 7982 58942 8034
rect 58942 7982 58994 8034
rect 58994 7982 58996 8034
rect 58940 7980 58996 7982
rect 59164 7644 59220 7700
rect 58604 6300 58660 6356
rect 58268 5964 58324 6020
rect 58604 5628 58660 5684
rect 58492 5234 58548 5236
rect 58492 5182 58494 5234
rect 58494 5182 58546 5234
rect 58546 5182 58548 5234
rect 58492 5180 58548 5182
rect 58940 4508 58996 4564
rect 57148 3442 57204 3444
rect 57148 3390 57150 3442
rect 57150 3390 57202 3442
rect 57202 3390 57204 3442
rect 57148 3388 57204 3390
rect 57036 2716 57092 2772
rect 58044 3388 58100 3444
rect 58940 3442 58996 3444
rect 58940 3390 58942 3442
rect 58942 3390 58994 3442
rect 58994 3390 58996 3442
rect 58940 3388 58996 3390
rect 58380 3276 58436 3332
rect 58380 2604 58436 2660
rect 59388 6578 59444 6580
rect 59388 6526 59390 6578
rect 59390 6526 59442 6578
rect 59442 6526 59444 6578
rect 59388 6524 59444 6526
rect 59724 7084 59780 7140
rect 59724 6636 59780 6692
rect 59612 5906 59668 5908
rect 59612 5854 59614 5906
rect 59614 5854 59666 5906
rect 59666 5854 59668 5906
rect 59612 5852 59668 5854
rect 59500 5180 59556 5236
rect 59724 4396 59780 4452
rect 60732 7532 60788 7588
rect 60956 7532 61012 7588
rect 60396 6466 60452 6468
rect 60396 6414 60398 6466
rect 60398 6414 60450 6466
rect 60450 6414 60452 6466
rect 60396 6412 60452 6414
rect 60396 6076 60452 6132
rect 60620 6188 60676 6244
rect 60844 6412 60900 6468
rect 60508 5964 60564 6020
rect 60620 4956 60676 5012
rect 60508 4450 60564 4452
rect 60508 4398 60510 4450
rect 60510 4398 60562 4450
rect 60562 4398 60564 4450
rect 60508 4396 60564 4398
rect 59724 3388 59780 3444
rect 61516 10780 61572 10836
rect 61068 6076 61124 6132
rect 61180 8988 61236 9044
rect 60956 4508 61012 4564
rect 61628 10610 61684 10612
rect 61628 10558 61630 10610
rect 61630 10558 61682 10610
rect 61682 10558 61684 10610
rect 61628 10556 61684 10558
rect 61964 11900 62020 11956
rect 63420 16268 63476 16324
rect 61628 9100 61684 9156
rect 62636 11004 62692 11060
rect 63196 11170 63252 11172
rect 63196 11118 63198 11170
rect 63198 11118 63250 11170
rect 63250 11118 63252 11170
rect 63196 11116 63252 11118
rect 61404 8258 61460 8260
rect 61404 8206 61406 8258
rect 61406 8206 61458 8258
rect 61458 8206 61460 8258
rect 61404 8204 61460 8206
rect 61292 7644 61348 7700
rect 61516 7980 61572 8036
rect 61404 7362 61460 7364
rect 61404 7310 61406 7362
rect 61406 7310 61458 7362
rect 61458 7310 61460 7362
rect 61404 7308 61460 7310
rect 61292 6018 61348 6020
rect 61292 5966 61294 6018
rect 61294 5966 61346 6018
rect 61346 5966 61348 6018
rect 61292 5964 61348 5966
rect 61852 6636 61908 6692
rect 61740 6466 61796 6468
rect 61740 6414 61742 6466
rect 61742 6414 61794 6466
rect 61794 6414 61796 6466
rect 61740 6412 61796 6414
rect 61628 6300 61684 6356
rect 61404 4844 61460 4900
rect 61852 5122 61908 5124
rect 61852 5070 61854 5122
rect 61854 5070 61906 5122
rect 61906 5070 61908 5122
rect 61852 5068 61908 5070
rect 60732 1484 60788 1540
rect 61852 4562 61908 4564
rect 61852 4510 61854 4562
rect 61854 4510 61906 4562
rect 61906 4510 61908 4562
rect 61852 4508 61908 4510
rect 62300 9884 62356 9940
rect 62636 10108 62692 10164
rect 62300 8988 62356 9044
rect 62524 9602 62580 9604
rect 62524 9550 62526 9602
rect 62526 9550 62578 9602
rect 62578 9550 62580 9602
rect 62524 9548 62580 9550
rect 62524 8988 62580 9044
rect 62188 8428 62244 8484
rect 62412 7698 62468 7700
rect 62412 7646 62414 7698
rect 62414 7646 62466 7698
rect 62466 7646 62468 7698
rect 62412 7644 62468 7646
rect 63756 12290 63812 12292
rect 63756 12238 63758 12290
rect 63758 12238 63810 12290
rect 63810 12238 63812 12290
rect 63756 12236 63812 12238
rect 63756 11506 63812 11508
rect 63756 11454 63758 11506
rect 63758 11454 63810 11506
rect 63810 11454 63812 11506
rect 63756 11452 63812 11454
rect 64540 12236 64596 12292
rect 63980 11340 64036 11396
rect 63196 10108 63252 10164
rect 63420 9938 63476 9940
rect 63420 9886 63422 9938
rect 63422 9886 63474 9938
rect 63474 9886 63476 9938
rect 63420 9884 63476 9886
rect 62972 9602 63028 9604
rect 62972 9550 62974 9602
rect 62974 9550 63026 9602
rect 63026 9550 63028 9602
rect 62972 9548 63028 9550
rect 63420 8988 63476 9044
rect 62860 8876 62916 8932
rect 62300 6636 62356 6692
rect 62972 6972 63028 7028
rect 62300 5346 62356 5348
rect 62300 5294 62302 5346
rect 62302 5294 62354 5346
rect 62354 5294 62356 5346
rect 62300 5292 62356 5294
rect 62636 6524 62692 6580
rect 62860 6300 62916 6356
rect 62748 5292 62804 5348
rect 62524 4956 62580 5012
rect 62076 4396 62132 4452
rect 62300 4620 62356 4676
rect 62860 5068 62916 5124
rect 63196 4844 63252 4900
rect 61516 3276 61572 3332
rect 62524 4284 62580 4340
rect 63980 10556 64036 10612
rect 63756 8428 63812 8484
rect 63868 9212 63924 9268
rect 64204 9212 64260 9268
rect 64204 8930 64260 8932
rect 64204 8878 64206 8930
rect 64206 8878 64258 8930
rect 64258 8878 64260 8930
rect 64204 8876 64260 8878
rect 63868 8092 63924 8148
rect 63532 6972 63588 7028
rect 63420 6636 63476 6692
rect 63420 6300 63476 6356
rect 63644 6018 63700 6020
rect 63644 5966 63646 6018
rect 63646 5966 63698 6018
rect 63698 5966 63700 6018
rect 63644 5964 63700 5966
rect 64428 9042 64484 9044
rect 64428 8990 64430 9042
rect 64430 8990 64482 9042
rect 64482 8990 64484 9042
rect 64428 8988 64484 8990
rect 64876 10668 64932 10724
rect 64764 10498 64820 10500
rect 64764 10446 64766 10498
rect 64766 10446 64818 10498
rect 64818 10446 64820 10498
rect 64764 10444 64820 10446
rect 64764 10108 64820 10164
rect 64652 8764 64708 8820
rect 64316 6412 64372 6468
rect 64092 6300 64148 6356
rect 64316 6188 64372 6244
rect 64428 5740 64484 5796
rect 64092 4844 64148 4900
rect 64316 4956 64372 5012
rect 64428 4732 64484 4788
rect 64428 4450 64484 4452
rect 64428 4398 64430 4450
rect 64430 4398 64482 4450
rect 64482 4398 64484 4450
rect 64428 4396 64484 4398
rect 63644 4060 63700 4116
rect 64652 4396 64708 4452
rect 64876 6636 64932 6692
rect 65436 12012 65492 12068
rect 65212 9548 65268 9604
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 67004 19292 67060 19348
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 66108 12066 66164 12068
rect 66108 12014 66110 12066
rect 66110 12014 66162 12066
rect 66162 12014 66164 12066
rect 66108 12012 66164 12014
rect 66892 12066 66948 12068
rect 66892 12014 66894 12066
rect 66894 12014 66946 12066
rect 66946 12014 66948 12066
rect 66892 12012 66948 12014
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 65660 11004 65716 11060
rect 66332 11004 66388 11060
rect 65548 10444 65604 10500
rect 65996 10668 66052 10724
rect 65916 10218 65972 10220
rect 65436 9602 65492 9604
rect 65436 9550 65438 9602
rect 65438 9550 65490 9602
rect 65490 9550 65492 9602
rect 65436 9548 65492 9550
rect 65548 10108 65604 10164
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 65436 9266 65492 9268
rect 65436 9214 65438 9266
rect 65438 9214 65490 9266
rect 65490 9214 65492 9266
rect 65436 9212 65492 9214
rect 65212 6188 65268 6244
rect 65324 9100 65380 9156
rect 65100 5964 65156 6020
rect 65100 5404 65156 5460
rect 64876 4172 64932 4228
rect 63532 3724 63588 3780
rect 64092 924 64148 980
rect 64764 3948 64820 4004
rect 64764 3666 64820 3668
rect 64764 3614 64766 3666
rect 64766 3614 64818 3666
rect 64818 3614 64820 3666
rect 64764 3612 64820 3614
rect 65772 9884 65828 9940
rect 66220 9266 66276 9268
rect 66220 9214 66222 9266
rect 66222 9214 66274 9266
rect 66274 9214 66276 9266
rect 66220 9212 66276 9214
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 66556 11116 66612 11172
rect 66556 9884 66612 9940
rect 66892 9266 66948 9268
rect 66892 9214 66894 9266
rect 66894 9214 66946 9266
rect 66946 9214 66948 9266
rect 66892 9212 66948 9214
rect 67116 11170 67172 11172
rect 67116 11118 67118 11170
rect 67118 11118 67170 11170
rect 67170 11118 67172 11170
rect 67116 11116 67172 11118
rect 67452 11004 67508 11060
rect 68796 25340 68852 25396
rect 68236 19740 68292 19796
rect 71372 116172 71428 116228
rect 69916 22652 69972 22708
rect 70140 28588 70196 28644
rect 69692 22092 69748 22148
rect 68796 13580 68852 13636
rect 69132 13634 69188 13636
rect 69132 13582 69134 13634
rect 69134 13582 69186 13634
rect 69186 13582 69188 13634
rect 69132 13580 69188 13582
rect 69580 13634 69636 13636
rect 69580 13582 69582 13634
rect 69582 13582 69634 13634
rect 69634 13582 69636 13634
rect 69580 13580 69636 13582
rect 67340 10668 67396 10724
rect 66444 8146 66500 8148
rect 66444 8094 66446 8146
rect 66446 8094 66498 8146
rect 66498 8094 66500 8146
rect 66444 8092 66500 8094
rect 66444 7420 66500 7476
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 65548 6130 65604 6132
rect 65548 6078 65550 6130
rect 65550 6078 65602 6130
rect 65602 6078 65604 6130
rect 65548 6076 65604 6078
rect 65660 6636 65716 6692
rect 65436 5794 65492 5796
rect 65436 5742 65438 5794
rect 65438 5742 65490 5794
rect 65490 5742 65492 5794
rect 65436 5740 65492 5742
rect 65548 5404 65604 5460
rect 65212 4620 65268 4676
rect 66108 6690 66164 6692
rect 66108 6638 66110 6690
rect 66110 6638 66162 6690
rect 66162 6638 66164 6690
rect 66108 6636 66164 6638
rect 65660 5180 65716 5236
rect 65772 6412 65828 6468
rect 66108 6188 66164 6244
rect 66556 6412 66612 6468
rect 66332 6018 66388 6020
rect 66332 5966 66334 6018
rect 66334 5966 66386 6018
rect 66386 5966 66388 6018
rect 66332 5964 66388 5966
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 66332 5292 66388 5348
rect 65772 4844 65828 4900
rect 66556 6188 66612 6244
rect 66444 4620 66500 4676
rect 66892 7474 66948 7476
rect 66892 7422 66894 7474
rect 66894 7422 66946 7474
rect 66946 7422 66948 7474
rect 66892 7420 66948 7422
rect 66668 5628 66724 5684
rect 66780 6524 66836 6580
rect 67004 6466 67060 6468
rect 67004 6414 67006 6466
rect 67006 6414 67058 6466
rect 67058 6414 67060 6466
rect 67004 6412 67060 6414
rect 66780 5740 66836 5796
rect 67564 10444 67620 10500
rect 67452 6300 67508 6356
rect 67228 6076 67284 6132
rect 68124 11170 68180 11172
rect 68124 11118 68126 11170
rect 68126 11118 68178 11170
rect 68178 11118 68180 11170
rect 68124 11116 68180 11118
rect 67788 10220 67844 10276
rect 67788 9266 67844 9268
rect 67788 9214 67790 9266
rect 67790 9214 67842 9266
rect 67842 9214 67844 9266
rect 67788 9212 67844 9214
rect 68124 10220 68180 10276
rect 67676 8876 67732 8932
rect 68460 12796 68516 12852
rect 68460 12348 68516 12404
rect 68348 9826 68404 9828
rect 68348 9774 68350 9826
rect 68350 9774 68402 9826
rect 68402 9774 68404 9826
rect 68348 9772 68404 9774
rect 68236 8652 68292 8708
rect 68012 7084 68068 7140
rect 67676 6578 67732 6580
rect 67676 6526 67678 6578
rect 67678 6526 67730 6578
rect 67730 6526 67732 6578
rect 67676 6524 67732 6526
rect 67788 6130 67844 6132
rect 67788 6078 67790 6130
rect 67790 6078 67842 6130
rect 67842 6078 67844 6130
rect 67788 6076 67844 6078
rect 67900 5964 67956 6020
rect 67564 5906 67620 5908
rect 67564 5854 67566 5906
rect 67566 5854 67618 5906
rect 67618 5854 67620 5906
rect 67564 5852 67620 5854
rect 67452 5628 67508 5684
rect 66668 4620 66724 4676
rect 67452 4844 67508 4900
rect 67676 5122 67732 5124
rect 67676 5070 67678 5122
rect 67678 5070 67730 5122
rect 67730 5070 67732 5122
rect 67676 5068 67732 5070
rect 67788 4844 67844 4900
rect 68124 6636 68180 6692
rect 68572 11340 68628 11396
rect 69132 11676 69188 11732
rect 68572 11170 68628 11172
rect 68572 11118 68574 11170
rect 68574 11118 68626 11170
rect 68626 11118 68628 11170
rect 68572 11116 68628 11118
rect 68684 11004 68740 11060
rect 68572 10892 68628 10948
rect 68572 9436 68628 9492
rect 68796 9772 68852 9828
rect 68684 9266 68740 9268
rect 68684 9214 68686 9266
rect 68686 9214 68738 9266
rect 68738 9214 68740 9266
rect 68684 9212 68740 9214
rect 68796 9436 68852 9492
rect 69020 8988 69076 9044
rect 68572 8930 68628 8932
rect 68572 8878 68574 8930
rect 68574 8878 68626 8930
rect 68626 8878 68628 8930
rect 68572 8876 68628 8878
rect 68796 8652 68852 8708
rect 69244 11170 69300 11172
rect 69244 11118 69246 11170
rect 69246 11118 69298 11170
rect 69298 11118 69300 11170
rect 69244 11116 69300 11118
rect 68908 7196 68964 7252
rect 69244 10556 69300 10612
rect 68796 6076 68852 6132
rect 68796 5628 68852 5684
rect 69692 11676 69748 11732
rect 69804 12012 69860 12068
rect 69692 11394 69748 11396
rect 69692 11342 69694 11394
rect 69694 11342 69746 11394
rect 69746 11342 69748 11394
rect 69692 11340 69748 11342
rect 72268 116226 72324 116228
rect 72268 116174 72270 116226
rect 72270 116174 72322 116226
rect 72322 116174 72324 116226
rect 72268 116172 72324 116174
rect 72604 115554 72660 115556
rect 72604 115502 72606 115554
rect 72606 115502 72658 115554
rect 72658 115502 72660 115554
rect 72604 115500 72660 115502
rect 71372 27356 71428 27412
rect 72156 25228 72212 25284
rect 70140 13074 70196 13076
rect 70140 13022 70142 13074
rect 70142 13022 70194 13074
rect 70194 13022 70196 13074
rect 70140 13020 70196 13022
rect 70252 23996 70308 24052
rect 71260 20524 71316 20580
rect 70252 12402 70308 12404
rect 70252 12350 70254 12402
rect 70254 12350 70306 12402
rect 70306 12350 70308 12402
rect 70252 12348 70308 12350
rect 70028 12012 70084 12068
rect 70588 12066 70644 12068
rect 70588 12014 70590 12066
rect 70590 12014 70642 12066
rect 70642 12014 70644 12066
rect 70588 12012 70644 12014
rect 71036 12908 71092 12964
rect 70924 12460 70980 12516
rect 70140 11506 70196 11508
rect 70140 11454 70142 11506
rect 70142 11454 70194 11506
rect 70194 11454 70196 11506
rect 70140 11452 70196 11454
rect 69692 8930 69748 8932
rect 69692 8878 69694 8930
rect 69694 8878 69746 8930
rect 69746 8878 69748 8930
rect 69692 8876 69748 8878
rect 70028 11340 70084 11396
rect 70028 8540 70084 8596
rect 69468 8092 69524 8148
rect 69356 7420 69412 7476
rect 69804 7308 69860 7364
rect 69692 7196 69748 7252
rect 69468 7084 69524 7140
rect 69356 6018 69412 6020
rect 69356 5966 69358 6018
rect 69358 5966 69410 6018
rect 69410 5966 69412 6018
rect 69356 5964 69412 5966
rect 68236 5234 68292 5236
rect 68236 5182 68238 5234
rect 68238 5182 68290 5234
rect 68290 5182 68292 5234
rect 68236 5180 68292 5182
rect 69580 5180 69636 5236
rect 68012 4844 68068 4900
rect 70028 6412 70084 6468
rect 70140 10892 70196 10948
rect 70812 11452 70868 11508
rect 70700 11394 70756 11396
rect 70700 11342 70702 11394
rect 70702 11342 70754 11394
rect 70754 11342 70756 11394
rect 70700 11340 70756 11342
rect 70252 10780 70308 10836
rect 70812 8540 70868 8596
rect 70252 5122 70308 5124
rect 70252 5070 70254 5122
rect 70254 5070 70306 5122
rect 70306 5070 70308 5122
rect 70252 5068 70308 5070
rect 70476 4956 70532 5012
rect 70588 6188 70644 6244
rect 70364 4844 70420 4900
rect 69356 4732 69412 4788
rect 68124 4620 68180 4676
rect 67900 4396 67956 4452
rect 68908 4620 68964 4676
rect 68348 4450 68404 4452
rect 68348 4398 68350 4450
rect 68350 4398 68402 4450
rect 68402 4398 68404 4450
rect 68348 4396 68404 4398
rect 69356 4338 69412 4340
rect 69356 4286 69358 4338
rect 69358 4286 69410 4338
rect 69410 4286 69412 4338
rect 69356 4284 69412 4286
rect 66108 4226 66164 4228
rect 66108 4174 66110 4226
rect 66110 4174 66162 4226
rect 66162 4174 66164 4226
rect 66108 4172 66164 4174
rect 69244 4172 69300 4228
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 66108 3724 66164 3780
rect 65548 3500 65604 3556
rect 68460 3554 68516 3556
rect 68460 3502 68462 3554
rect 68462 3502 68514 3554
rect 68514 3502 68516 3554
rect 68460 3500 68516 3502
rect 65884 3388 65940 3444
rect 64652 1036 64708 1092
rect 67004 3442 67060 3444
rect 67004 3390 67006 3442
rect 67006 3390 67058 3442
rect 67058 3390 67060 3442
rect 67004 3388 67060 3390
rect 67564 3388 67620 3444
rect 70028 4226 70084 4228
rect 70028 4174 70030 4226
rect 70030 4174 70082 4226
rect 70082 4174 70084 4226
rect 70028 4172 70084 4174
rect 70588 4732 70644 4788
rect 70700 5852 70756 5908
rect 69356 3442 69412 3444
rect 69356 3390 69358 3442
rect 69358 3390 69410 3442
rect 69410 3390 69412 3442
rect 69356 3388 69412 3390
rect 71036 12066 71092 12068
rect 71036 12014 71038 12066
rect 71038 12014 71090 12066
rect 71090 12014 71092 12066
rect 71036 12012 71092 12014
rect 71036 11788 71092 11844
rect 71260 10892 71316 10948
rect 71372 13580 71428 13636
rect 71036 7308 71092 7364
rect 71148 10332 71204 10388
rect 70924 6412 70980 6468
rect 70812 4844 70868 4900
rect 71036 5010 71092 5012
rect 71036 4958 71038 5010
rect 71038 4958 71090 5010
rect 71090 4958 71092 5010
rect 71036 4956 71092 4958
rect 70924 4396 70980 4452
rect 71260 9996 71316 10052
rect 71260 8092 71316 8148
rect 71260 7420 71316 7476
rect 71260 6972 71316 7028
rect 72940 15260 72996 15316
rect 72716 13634 72772 13636
rect 72716 13582 72718 13634
rect 72718 13582 72770 13634
rect 72770 13582 72772 13634
rect 72716 13580 72772 13582
rect 71484 12908 71540 12964
rect 71596 11676 71652 11732
rect 72156 12460 72212 12516
rect 72268 12348 72324 12404
rect 71932 11676 71988 11732
rect 71708 11340 71764 11396
rect 71596 11170 71652 11172
rect 71596 11118 71598 11170
rect 71598 11118 71650 11170
rect 71650 11118 71652 11170
rect 71596 11116 71652 11118
rect 71484 10780 71540 10836
rect 71820 10108 71876 10164
rect 71932 9996 71988 10052
rect 71596 7474 71652 7476
rect 71596 7422 71598 7474
rect 71598 7422 71650 7474
rect 71650 7422 71652 7474
rect 71596 7420 71652 7422
rect 71708 7362 71764 7364
rect 71708 7310 71710 7362
rect 71710 7310 71762 7362
rect 71762 7310 71764 7362
rect 71708 7308 71764 7310
rect 71932 6188 71988 6244
rect 72044 6412 72100 6468
rect 71372 5628 71428 5684
rect 71932 5292 71988 5348
rect 71260 5010 71316 5012
rect 71260 4958 71262 5010
rect 71262 4958 71314 5010
rect 71314 4958 71316 5010
rect 71260 4956 71316 4958
rect 71708 5180 71764 5236
rect 71372 4562 71428 4564
rect 71372 4510 71374 4562
rect 71374 4510 71426 4562
rect 71426 4510 71428 4562
rect 71372 4508 71428 4510
rect 71820 4450 71876 4452
rect 71820 4398 71822 4450
rect 71822 4398 71874 4450
rect 71874 4398 71876 4450
rect 71820 4396 71876 4398
rect 72716 9324 72772 9380
rect 72492 9042 72548 9044
rect 72492 8990 72494 9042
rect 72494 8990 72546 9042
rect 72546 8990 72548 9042
rect 72492 8988 72548 8990
rect 72268 8876 72324 8932
rect 72268 6076 72324 6132
rect 72380 5964 72436 6020
rect 72492 4844 72548 4900
rect 72604 4396 72660 4452
rect 72380 4338 72436 4340
rect 72380 4286 72382 4338
rect 72382 4286 72434 4338
rect 72434 4286 72436 4338
rect 72380 4284 72436 4286
rect 73500 116508 73556 116564
rect 74396 116562 74452 116564
rect 74396 116510 74398 116562
rect 74398 116510 74450 116562
rect 74450 116510 74452 116562
rect 74396 116508 74452 116510
rect 75068 116508 75124 116564
rect 76524 116562 76580 116564
rect 76524 116510 76526 116562
rect 76526 116510 76578 116562
rect 76578 116510 76580 116562
rect 76524 116508 76580 116510
rect 78204 116620 78260 116676
rect 78988 116620 79044 116676
rect 79772 116508 79828 116564
rect 80668 116562 80724 116564
rect 80668 116510 80670 116562
rect 80670 116510 80722 116562
rect 80722 116510 80724 116562
rect 80668 116508 80724 116510
rect 73500 115500 73556 115556
rect 77308 115554 77364 115556
rect 77308 115502 77310 115554
rect 77310 115502 77362 115554
rect 77362 115502 77364 115554
rect 77308 115500 77364 115502
rect 77980 115500 78036 115556
rect 74844 29372 74900 29428
rect 74732 22428 74788 22484
rect 73948 22204 74004 22260
rect 73948 13468 74004 13524
rect 74060 14364 74116 14420
rect 73052 12012 73108 12068
rect 73612 12290 73668 12292
rect 73612 12238 73614 12290
rect 73614 12238 73666 12290
rect 73666 12238 73668 12290
rect 73612 12236 73668 12238
rect 73276 11116 73332 11172
rect 73500 11116 73556 11172
rect 73388 10610 73444 10612
rect 73388 10558 73390 10610
rect 73390 10558 73442 10610
rect 73442 10558 73444 10610
rect 73388 10556 73444 10558
rect 73164 5852 73220 5908
rect 73276 9324 73332 9380
rect 72940 4284 72996 4340
rect 73836 10780 73892 10836
rect 73724 10668 73780 10724
rect 73836 10444 73892 10500
rect 73724 9266 73780 9268
rect 73724 9214 73726 9266
rect 73726 9214 73778 9266
rect 73778 9214 73780 9266
rect 73724 9212 73780 9214
rect 74956 22316 75012 22372
rect 76076 20972 76132 21028
rect 74844 13020 74900 13076
rect 74172 12348 74228 12404
rect 74172 11452 74228 11508
rect 74172 10668 74228 10724
rect 74060 8988 74116 9044
rect 73836 8428 73892 8484
rect 74060 6018 74116 6020
rect 74060 5966 74062 6018
rect 74062 5966 74114 6018
rect 74114 5966 74116 6018
rect 74060 5964 74116 5966
rect 73388 5906 73444 5908
rect 73388 5854 73390 5906
rect 73390 5854 73442 5906
rect 73442 5854 73444 5906
rect 73388 5852 73444 5854
rect 73948 5906 74004 5908
rect 73948 5854 73950 5906
rect 73950 5854 74002 5906
rect 74002 5854 74004 5906
rect 73948 5852 74004 5854
rect 73500 5068 73556 5124
rect 73612 4956 73668 5012
rect 73612 4508 73668 4564
rect 70700 1148 70756 1204
rect 73836 5068 73892 5124
rect 73612 3612 73668 3668
rect 74060 4450 74116 4452
rect 74060 4398 74062 4450
rect 74062 4398 74114 4450
rect 74114 4398 74116 4450
rect 74060 4396 74116 4398
rect 74956 12460 75012 12516
rect 74508 11788 74564 11844
rect 74956 10722 75012 10724
rect 74956 10670 74958 10722
rect 74958 10670 75010 10722
rect 75010 10670 75012 10722
rect 74956 10668 75012 10670
rect 74844 10610 74900 10612
rect 74844 10558 74846 10610
rect 74846 10558 74898 10610
rect 74898 10558 74900 10610
rect 74844 10556 74900 10558
rect 74732 9660 74788 9716
rect 74620 8988 74676 9044
rect 74508 8204 74564 8260
rect 74508 7474 74564 7476
rect 74508 7422 74510 7474
rect 74510 7422 74562 7474
rect 74562 7422 74564 7474
rect 74508 7420 74564 7422
rect 74732 5794 74788 5796
rect 74732 5742 74734 5794
rect 74734 5742 74786 5794
rect 74786 5742 74788 5794
rect 74732 5740 74788 5742
rect 74396 4338 74452 4340
rect 74396 4286 74398 4338
rect 74398 4286 74450 4338
rect 74450 4286 74452 4338
rect 74396 4284 74452 4286
rect 74620 4060 74676 4116
rect 74396 3388 74452 3444
rect 74620 2604 74676 2660
rect 75404 13468 75460 13524
rect 75628 13468 75684 13524
rect 75180 12738 75236 12740
rect 75180 12686 75182 12738
rect 75182 12686 75234 12738
rect 75234 12686 75236 12738
rect 75180 12684 75236 12686
rect 75292 10108 75348 10164
rect 75180 9714 75236 9716
rect 75180 9662 75182 9714
rect 75182 9662 75234 9714
rect 75234 9662 75236 9714
rect 75180 9660 75236 9662
rect 75292 9436 75348 9492
rect 75404 9212 75460 9268
rect 75404 9042 75460 9044
rect 75404 8990 75406 9042
rect 75406 8990 75458 9042
rect 75458 8990 75460 9042
rect 75404 8988 75460 8990
rect 75964 12796 76020 12852
rect 75852 12348 75908 12404
rect 75404 8428 75460 8484
rect 75292 8316 75348 8372
rect 75516 8316 75572 8372
rect 75516 7756 75572 7812
rect 75404 7698 75460 7700
rect 75404 7646 75406 7698
rect 75406 7646 75458 7698
rect 75458 7646 75460 7698
rect 75404 7644 75460 7646
rect 75516 7532 75572 7588
rect 75292 7474 75348 7476
rect 75292 7422 75294 7474
rect 75294 7422 75346 7474
rect 75346 7422 75348 7474
rect 75292 7420 75348 7422
rect 75292 7196 75348 7252
rect 75068 5404 75124 5460
rect 75740 12012 75796 12068
rect 75740 11340 75796 11396
rect 77868 20748 77924 20804
rect 77644 15820 77700 15876
rect 77308 13804 77364 13860
rect 77084 13634 77140 13636
rect 77084 13582 77086 13634
rect 77086 13582 77138 13634
rect 77138 13582 77140 13634
rect 77084 13580 77140 13582
rect 76076 12402 76132 12404
rect 76076 12350 76078 12402
rect 76078 12350 76130 12402
rect 76130 12350 76132 12402
rect 76076 12348 76132 12350
rect 76188 12572 76244 12628
rect 76188 12124 76244 12180
rect 76188 11004 76244 11060
rect 76188 10668 76244 10724
rect 76188 10498 76244 10500
rect 76188 10446 76190 10498
rect 76190 10446 76242 10498
rect 76242 10446 76244 10498
rect 76188 10444 76244 10446
rect 76300 9212 76356 9268
rect 77084 13132 77140 13188
rect 77196 13468 77252 13524
rect 76524 13020 76580 13076
rect 76636 12962 76692 12964
rect 76636 12910 76638 12962
rect 76638 12910 76690 12962
rect 76690 12910 76692 12962
rect 76636 12908 76692 12910
rect 77084 12796 77140 12852
rect 77084 12402 77140 12404
rect 77084 12350 77086 12402
rect 77086 12350 77138 12402
rect 77138 12350 77140 12402
rect 77084 12348 77140 12350
rect 77196 12236 77252 12292
rect 75852 8316 75908 8372
rect 75740 7756 75796 7812
rect 75628 7196 75684 7252
rect 75404 6076 75460 6132
rect 76524 8146 76580 8148
rect 76524 8094 76526 8146
rect 76526 8094 76578 8146
rect 76578 8094 76580 8146
rect 76524 8092 76580 8094
rect 75964 6524 76020 6580
rect 76524 7756 76580 7812
rect 75516 5852 75572 5908
rect 75404 5292 75460 5348
rect 75292 5234 75348 5236
rect 75292 5182 75294 5234
rect 75294 5182 75346 5234
rect 75346 5182 75348 5234
rect 75292 5180 75348 5182
rect 75180 5068 75236 5124
rect 74956 4284 75012 4340
rect 75628 5292 75684 5348
rect 75516 5068 75572 5124
rect 76524 7308 76580 7364
rect 76188 6748 76244 6804
rect 76412 6972 76468 7028
rect 76636 6636 76692 6692
rect 76524 6524 76580 6580
rect 76188 5180 76244 5236
rect 76860 9436 76916 9492
rect 76972 12012 77028 12068
rect 77196 11506 77252 11508
rect 77196 11454 77198 11506
rect 77198 11454 77250 11506
rect 77250 11454 77252 11506
rect 77196 11452 77252 11454
rect 77196 9772 77252 9828
rect 77084 7308 77140 7364
rect 77420 13020 77476 13076
rect 77420 12012 77476 12068
rect 80220 116060 80276 116116
rect 78876 23884 78932 23940
rect 78204 18508 78260 18564
rect 77532 11452 77588 11508
rect 77532 9212 77588 9268
rect 77420 8764 77476 8820
rect 77756 9826 77812 9828
rect 77756 9774 77758 9826
rect 77758 9774 77810 9826
rect 77810 9774 77812 9826
rect 77756 9772 77812 9774
rect 77980 12402 78036 12404
rect 77980 12350 77982 12402
rect 77982 12350 78034 12402
rect 78034 12350 78036 12402
rect 77980 12348 78036 12350
rect 79436 23548 79492 23604
rect 78876 13580 78932 13636
rect 79100 13634 79156 13636
rect 79100 13582 79102 13634
rect 79102 13582 79154 13634
rect 79154 13582 79156 13634
rect 79100 13580 79156 13582
rect 78764 13468 78820 13524
rect 78540 12460 78596 12516
rect 78316 11788 78372 11844
rect 78092 11506 78148 11508
rect 78092 11454 78094 11506
rect 78094 11454 78146 11506
rect 78146 11454 78148 11506
rect 78092 11452 78148 11454
rect 78204 11340 78260 11396
rect 78204 8930 78260 8932
rect 78204 8878 78206 8930
rect 78206 8878 78258 8930
rect 78258 8878 78260 8930
rect 78204 8876 78260 8878
rect 79436 12684 79492 12740
rect 79100 11788 79156 11844
rect 79212 12124 79268 12180
rect 78540 11452 78596 11508
rect 78428 11394 78484 11396
rect 78428 11342 78430 11394
rect 78430 11342 78482 11394
rect 78482 11342 78484 11394
rect 78428 11340 78484 11342
rect 78316 11004 78372 11060
rect 78876 10444 78932 10500
rect 78428 10220 78484 10276
rect 79324 11452 79380 11508
rect 78764 9714 78820 9716
rect 78764 9662 78766 9714
rect 78766 9662 78818 9714
rect 78818 9662 78820 9714
rect 78764 9660 78820 9662
rect 79212 9714 79268 9716
rect 79212 9662 79214 9714
rect 79214 9662 79266 9714
rect 79266 9662 79268 9714
rect 79212 9660 79268 9662
rect 78540 9212 78596 9268
rect 78428 9100 78484 9156
rect 78764 8930 78820 8932
rect 78764 8878 78766 8930
rect 78766 8878 78818 8930
rect 78818 8878 78820 8930
rect 78764 8876 78820 8878
rect 78316 8652 78372 8708
rect 77532 7868 77588 7924
rect 77756 7756 77812 7812
rect 77644 7420 77700 7476
rect 77308 6860 77364 6916
rect 77532 7196 77588 7252
rect 77532 6802 77588 6804
rect 77532 6750 77534 6802
rect 77534 6750 77586 6802
rect 77586 6750 77588 6802
rect 77532 6748 77588 6750
rect 77308 6690 77364 6692
rect 77308 6638 77310 6690
rect 77310 6638 77362 6690
rect 77362 6638 77364 6690
rect 77308 6636 77364 6638
rect 77420 6466 77476 6468
rect 77420 6414 77422 6466
rect 77422 6414 77474 6466
rect 77474 6414 77476 6466
rect 77420 6412 77476 6414
rect 77756 6524 77812 6580
rect 77756 6188 77812 6244
rect 76972 5292 77028 5348
rect 77644 5122 77700 5124
rect 77644 5070 77646 5122
rect 77646 5070 77698 5122
rect 77698 5070 77700 5122
rect 77644 5068 77700 5070
rect 77084 4956 77140 5012
rect 76748 4844 76804 4900
rect 76524 4732 76580 4788
rect 77308 4732 77364 4788
rect 76300 4172 76356 4228
rect 76300 3948 76356 4004
rect 76524 4508 76580 4564
rect 74844 3836 74900 3892
rect 75964 3724 76020 3780
rect 75180 3442 75236 3444
rect 75180 3390 75182 3442
rect 75182 3390 75234 3442
rect 75234 3390 75236 3442
rect 75180 3388 75236 3390
rect 74732 2492 74788 2548
rect 76860 3724 76916 3780
rect 76972 3836 77028 3892
rect 77084 3666 77140 3668
rect 77084 3614 77086 3666
rect 77086 3614 77138 3666
rect 77138 3614 77140 3666
rect 77084 3612 77140 3614
rect 77420 4620 77476 4676
rect 77532 3612 77588 3668
rect 78204 7196 78260 7252
rect 78540 8370 78596 8372
rect 78540 8318 78542 8370
rect 78542 8318 78594 8370
rect 78594 8318 78596 8370
rect 78540 8316 78596 8318
rect 78428 7756 78484 7812
rect 78540 8092 78596 8148
rect 78988 8258 79044 8260
rect 78988 8206 78990 8258
rect 78990 8206 79042 8258
rect 79042 8206 79044 8258
rect 78988 8204 79044 8206
rect 78876 7868 78932 7924
rect 78092 6860 78148 6916
rect 77980 6300 78036 6356
rect 77980 5906 78036 5908
rect 77980 5854 77982 5906
rect 77982 5854 78034 5906
rect 78034 5854 78036 5906
rect 77980 5852 78036 5854
rect 78428 6578 78484 6580
rect 78428 6526 78430 6578
rect 78430 6526 78482 6578
rect 78482 6526 78484 6578
rect 78428 6524 78484 6526
rect 77980 5010 78036 5012
rect 77980 4958 77982 5010
rect 77982 4958 78034 5010
rect 78034 4958 78036 5010
rect 77980 4956 78036 4958
rect 78092 4898 78148 4900
rect 78092 4846 78094 4898
rect 78094 4846 78146 4898
rect 78146 4846 78148 4898
rect 78092 4844 78148 4846
rect 78204 4396 78260 4452
rect 78428 4844 78484 4900
rect 79212 7868 79268 7924
rect 78876 6188 78932 6244
rect 78988 5852 79044 5908
rect 78652 5234 78708 5236
rect 78652 5182 78654 5234
rect 78654 5182 78706 5234
rect 78706 5182 78708 5234
rect 78652 5180 78708 5182
rect 78652 4956 78708 5012
rect 78652 4732 78708 4788
rect 79436 6860 79492 6916
rect 80780 22988 80836 23044
rect 80220 13468 80276 13524
rect 80556 16828 80612 16884
rect 79660 12850 79716 12852
rect 79660 12798 79662 12850
rect 79662 12798 79714 12850
rect 79714 12798 79716 12850
rect 79660 12796 79716 12798
rect 79884 12796 79940 12852
rect 79660 11788 79716 11844
rect 79772 10444 79828 10500
rect 79660 9436 79716 9492
rect 79660 9266 79716 9268
rect 79660 9214 79662 9266
rect 79662 9214 79714 9266
rect 79714 9214 79716 9266
rect 79660 9212 79716 9214
rect 79996 12460 80052 12516
rect 79772 7644 79828 7700
rect 79884 8146 79940 8148
rect 79884 8094 79886 8146
rect 79886 8094 79938 8146
rect 79938 8094 79940 8146
rect 79884 8092 79940 8094
rect 79884 7532 79940 7588
rect 79772 6860 79828 6916
rect 80108 12066 80164 12068
rect 80108 12014 80110 12066
rect 80110 12014 80162 12066
rect 80162 12014 80164 12066
rect 80108 12012 80164 12014
rect 80108 9602 80164 9604
rect 80108 9550 80110 9602
rect 80110 9550 80162 9602
rect 80162 9550 80164 9602
rect 80108 9548 80164 9550
rect 80108 8930 80164 8932
rect 80108 8878 80110 8930
rect 80110 8878 80162 8930
rect 80162 8878 80164 8930
rect 80108 8876 80164 8878
rect 80108 8540 80164 8596
rect 79772 6578 79828 6580
rect 79772 6526 79774 6578
rect 79774 6526 79826 6578
rect 79826 6526 79828 6578
rect 79772 6524 79828 6526
rect 79884 6300 79940 6356
rect 80108 6076 80164 6132
rect 79996 5964 80052 6020
rect 80556 12460 80612 12516
rect 80444 9212 80500 9268
rect 80444 8428 80500 8484
rect 80556 8764 80612 8820
rect 81276 116058 81332 116060
rect 81276 116006 81278 116058
rect 81278 116006 81330 116058
rect 81330 116006 81332 116058
rect 81276 116004 81332 116006
rect 81380 116058 81436 116060
rect 81380 116006 81382 116058
rect 81382 116006 81434 116058
rect 81434 116006 81436 116058
rect 81380 116004 81436 116006
rect 81484 116058 81540 116060
rect 81484 116006 81486 116058
rect 81486 116006 81538 116058
rect 81538 116006 81540 116058
rect 81484 116004 81540 116006
rect 85932 116060 85988 116116
rect 86380 116060 86436 116116
rect 82908 115836 82964 115892
rect 83804 115836 83860 115892
rect 81676 115554 81732 115556
rect 81676 115502 81678 115554
rect 81678 115502 81730 115554
rect 81730 115502 81732 115554
rect 81676 115500 81732 115502
rect 82236 115500 82292 115556
rect 82236 114828 82292 114884
rect 86716 114882 86772 114884
rect 86716 114830 86718 114882
rect 86718 114830 86770 114882
rect 86770 114830 86772 114882
rect 86716 114828 86772 114830
rect 92316 116620 92372 116676
rect 93212 116620 93268 116676
rect 90636 116172 90692 116228
rect 91084 116226 91140 116228
rect 91084 116174 91086 116226
rect 91086 116174 91138 116226
rect 91138 116174 91140 116226
rect 91084 116172 91140 116174
rect 90860 116060 90916 116116
rect 87612 114882 87668 114884
rect 87612 114830 87614 114882
rect 87614 114830 87666 114882
rect 87666 114830 87668 114882
rect 87612 114828 87668 114830
rect 81276 114490 81332 114492
rect 81276 114438 81278 114490
rect 81278 114438 81330 114490
rect 81330 114438 81332 114490
rect 81276 114436 81332 114438
rect 81380 114490 81436 114492
rect 81380 114438 81382 114490
rect 81382 114438 81434 114490
rect 81434 114438 81436 114490
rect 81380 114436 81436 114438
rect 81484 114490 81540 114492
rect 81484 114438 81486 114490
rect 81486 114438 81538 114490
rect 81538 114438 81540 114490
rect 81484 114436 81540 114438
rect 81276 112922 81332 112924
rect 81276 112870 81278 112922
rect 81278 112870 81330 112922
rect 81330 112870 81332 112922
rect 81276 112868 81332 112870
rect 81380 112922 81436 112924
rect 81380 112870 81382 112922
rect 81382 112870 81434 112922
rect 81434 112870 81436 112922
rect 81380 112868 81436 112870
rect 81484 112922 81540 112924
rect 81484 112870 81486 112922
rect 81486 112870 81538 112922
rect 81538 112870 81540 112922
rect 81484 112868 81540 112870
rect 81276 111354 81332 111356
rect 81276 111302 81278 111354
rect 81278 111302 81330 111354
rect 81330 111302 81332 111354
rect 81276 111300 81332 111302
rect 81380 111354 81436 111356
rect 81380 111302 81382 111354
rect 81382 111302 81434 111354
rect 81434 111302 81436 111354
rect 81380 111300 81436 111302
rect 81484 111354 81540 111356
rect 81484 111302 81486 111354
rect 81486 111302 81538 111354
rect 81538 111302 81540 111354
rect 81484 111300 81540 111302
rect 81276 109786 81332 109788
rect 81276 109734 81278 109786
rect 81278 109734 81330 109786
rect 81330 109734 81332 109786
rect 81276 109732 81332 109734
rect 81380 109786 81436 109788
rect 81380 109734 81382 109786
rect 81382 109734 81434 109786
rect 81434 109734 81436 109786
rect 81380 109732 81436 109734
rect 81484 109786 81540 109788
rect 81484 109734 81486 109786
rect 81486 109734 81538 109786
rect 81538 109734 81540 109786
rect 81484 109732 81540 109734
rect 81276 108218 81332 108220
rect 81276 108166 81278 108218
rect 81278 108166 81330 108218
rect 81330 108166 81332 108218
rect 81276 108164 81332 108166
rect 81380 108218 81436 108220
rect 81380 108166 81382 108218
rect 81382 108166 81434 108218
rect 81434 108166 81436 108218
rect 81380 108164 81436 108166
rect 81484 108218 81540 108220
rect 81484 108166 81486 108218
rect 81486 108166 81538 108218
rect 81538 108166 81540 108218
rect 81484 108164 81540 108166
rect 81276 106650 81332 106652
rect 81276 106598 81278 106650
rect 81278 106598 81330 106650
rect 81330 106598 81332 106650
rect 81276 106596 81332 106598
rect 81380 106650 81436 106652
rect 81380 106598 81382 106650
rect 81382 106598 81434 106650
rect 81434 106598 81436 106650
rect 81380 106596 81436 106598
rect 81484 106650 81540 106652
rect 81484 106598 81486 106650
rect 81486 106598 81538 106650
rect 81538 106598 81540 106650
rect 81484 106596 81540 106598
rect 81276 105082 81332 105084
rect 81276 105030 81278 105082
rect 81278 105030 81330 105082
rect 81330 105030 81332 105082
rect 81276 105028 81332 105030
rect 81380 105082 81436 105084
rect 81380 105030 81382 105082
rect 81382 105030 81434 105082
rect 81434 105030 81436 105082
rect 81380 105028 81436 105030
rect 81484 105082 81540 105084
rect 81484 105030 81486 105082
rect 81486 105030 81538 105082
rect 81538 105030 81540 105082
rect 81484 105028 81540 105030
rect 81276 103514 81332 103516
rect 81276 103462 81278 103514
rect 81278 103462 81330 103514
rect 81330 103462 81332 103514
rect 81276 103460 81332 103462
rect 81380 103514 81436 103516
rect 81380 103462 81382 103514
rect 81382 103462 81434 103514
rect 81434 103462 81436 103514
rect 81380 103460 81436 103462
rect 81484 103514 81540 103516
rect 81484 103462 81486 103514
rect 81486 103462 81538 103514
rect 81538 103462 81540 103514
rect 81484 103460 81540 103462
rect 81276 101946 81332 101948
rect 81276 101894 81278 101946
rect 81278 101894 81330 101946
rect 81330 101894 81332 101946
rect 81276 101892 81332 101894
rect 81380 101946 81436 101948
rect 81380 101894 81382 101946
rect 81382 101894 81434 101946
rect 81434 101894 81436 101946
rect 81380 101892 81436 101894
rect 81484 101946 81540 101948
rect 81484 101894 81486 101946
rect 81486 101894 81538 101946
rect 81538 101894 81540 101946
rect 81484 101892 81540 101894
rect 81276 100378 81332 100380
rect 81276 100326 81278 100378
rect 81278 100326 81330 100378
rect 81330 100326 81332 100378
rect 81276 100324 81332 100326
rect 81380 100378 81436 100380
rect 81380 100326 81382 100378
rect 81382 100326 81434 100378
rect 81434 100326 81436 100378
rect 81380 100324 81436 100326
rect 81484 100378 81540 100380
rect 81484 100326 81486 100378
rect 81486 100326 81538 100378
rect 81538 100326 81540 100378
rect 81484 100324 81540 100326
rect 81276 98810 81332 98812
rect 81276 98758 81278 98810
rect 81278 98758 81330 98810
rect 81330 98758 81332 98810
rect 81276 98756 81332 98758
rect 81380 98810 81436 98812
rect 81380 98758 81382 98810
rect 81382 98758 81434 98810
rect 81434 98758 81436 98810
rect 81380 98756 81436 98758
rect 81484 98810 81540 98812
rect 81484 98758 81486 98810
rect 81486 98758 81538 98810
rect 81538 98758 81540 98810
rect 81484 98756 81540 98758
rect 81276 97242 81332 97244
rect 81276 97190 81278 97242
rect 81278 97190 81330 97242
rect 81330 97190 81332 97242
rect 81276 97188 81332 97190
rect 81380 97242 81436 97244
rect 81380 97190 81382 97242
rect 81382 97190 81434 97242
rect 81434 97190 81436 97242
rect 81380 97188 81436 97190
rect 81484 97242 81540 97244
rect 81484 97190 81486 97242
rect 81486 97190 81538 97242
rect 81538 97190 81540 97242
rect 81484 97188 81540 97190
rect 81276 95674 81332 95676
rect 81276 95622 81278 95674
rect 81278 95622 81330 95674
rect 81330 95622 81332 95674
rect 81276 95620 81332 95622
rect 81380 95674 81436 95676
rect 81380 95622 81382 95674
rect 81382 95622 81434 95674
rect 81434 95622 81436 95674
rect 81380 95620 81436 95622
rect 81484 95674 81540 95676
rect 81484 95622 81486 95674
rect 81486 95622 81538 95674
rect 81538 95622 81540 95674
rect 81484 95620 81540 95622
rect 81276 94106 81332 94108
rect 81276 94054 81278 94106
rect 81278 94054 81330 94106
rect 81330 94054 81332 94106
rect 81276 94052 81332 94054
rect 81380 94106 81436 94108
rect 81380 94054 81382 94106
rect 81382 94054 81434 94106
rect 81434 94054 81436 94106
rect 81380 94052 81436 94054
rect 81484 94106 81540 94108
rect 81484 94054 81486 94106
rect 81486 94054 81538 94106
rect 81538 94054 81540 94106
rect 81484 94052 81540 94054
rect 81276 92538 81332 92540
rect 81276 92486 81278 92538
rect 81278 92486 81330 92538
rect 81330 92486 81332 92538
rect 81276 92484 81332 92486
rect 81380 92538 81436 92540
rect 81380 92486 81382 92538
rect 81382 92486 81434 92538
rect 81434 92486 81436 92538
rect 81380 92484 81436 92486
rect 81484 92538 81540 92540
rect 81484 92486 81486 92538
rect 81486 92486 81538 92538
rect 81538 92486 81540 92538
rect 81484 92484 81540 92486
rect 81276 90970 81332 90972
rect 81276 90918 81278 90970
rect 81278 90918 81330 90970
rect 81330 90918 81332 90970
rect 81276 90916 81332 90918
rect 81380 90970 81436 90972
rect 81380 90918 81382 90970
rect 81382 90918 81434 90970
rect 81434 90918 81436 90970
rect 81380 90916 81436 90918
rect 81484 90970 81540 90972
rect 81484 90918 81486 90970
rect 81486 90918 81538 90970
rect 81538 90918 81540 90970
rect 81484 90916 81540 90918
rect 81276 89402 81332 89404
rect 81276 89350 81278 89402
rect 81278 89350 81330 89402
rect 81330 89350 81332 89402
rect 81276 89348 81332 89350
rect 81380 89402 81436 89404
rect 81380 89350 81382 89402
rect 81382 89350 81434 89402
rect 81434 89350 81436 89402
rect 81380 89348 81436 89350
rect 81484 89402 81540 89404
rect 81484 89350 81486 89402
rect 81486 89350 81538 89402
rect 81538 89350 81540 89402
rect 81484 89348 81540 89350
rect 81276 87834 81332 87836
rect 81276 87782 81278 87834
rect 81278 87782 81330 87834
rect 81330 87782 81332 87834
rect 81276 87780 81332 87782
rect 81380 87834 81436 87836
rect 81380 87782 81382 87834
rect 81382 87782 81434 87834
rect 81434 87782 81436 87834
rect 81380 87780 81436 87782
rect 81484 87834 81540 87836
rect 81484 87782 81486 87834
rect 81486 87782 81538 87834
rect 81538 87782 81540 87834
rect 81484 87780 81540 87782
rect 81276 86266 81332 86268
rect 81276 86214 81278 86266
rect 81278 86214 81330 86266
rect 81330 86214 81332 86266
rect 81276 86212 81332 86214
rect 81380 86266 81436 86268
rect 81380 86214 81382 86266
rect 81382 86214 81434 86266
rect 81434 86214 81436 86266
rect 81380 86212 81436 86214
rect 81484 86266 81540 86268
rect 81484 86214 81486 86266
rect 81486 86214 81538 86266
rect 81538 86214 81540 86266
rect 81484 86212 81540 86214
rect 81276 84698 81332 84700
rect 81276 84646 81278 84698
rect 81278 84646 81330 84698
rect 81330 84646 81332 84698
rect 81276 84644 81332 84646
rect 81380 84698 81436 84700
rect 81380 84646 81382 84698
rect 81382 84646 81434 84698
rect 81434 84646 81436 84698
rect 81380 84644 81436 84646
rect 81484 84698 81540 84700
rect 81484 84646 81486 84698
rect 81486 84646 81538 84698
rect 81538 84646 81540 84698
rect 81484 84644 81540 84646
rect 81276 83130 81332 83132
rect 81276 83078 81278 83130
rect 81278 83078 81330 83130
rect 81330 83078 81332 83130
rect 81276 83076 81332 83078
rect 81380 83130 81436 83132
rect 81380 83078 81382 83130
rect 81382 83078 81434 83130
rect 81434 83078 81436 83130
rect 81380 83076 81436 83078
rect 81484 83130 81540 83132
rect 81484 83078 81486 83130
rect 81486 83078 81538 83130
rect 81538 83078 81540 83130
rect 81484 83076 81540 83078
rect 81276 81562 81332 81564
rect 81276 81510 81278 81562
rect 81278 81510 81330 81562
rect 81330 81510 81332 81562
rect 81276 81508 81332 81510
rect 81380 81562 81436 81564
rect 81380 81510 81382 81562
rect 81382 81510 81434 81562
rect 81434 81510 81436 81562
rect 81380 81508 81436 81510
rect 81484 81562 81540 81564
rect 81484 81510 81486 81562
rect 81486 81510 81538 81562
rect 81538 81510 81540 81562
rect 81484 81508 81540 81510
rect 81276 79994 81332 79996
rect 81276 79942 81278 79994
rect 81278 79942 81330 79994
rect 81330 79942 81332 79994
rect 81276 79940 81332 79942
rect 81380 79994 81436 79996
rect 81380 79942 81382 79994
rect 81382 79942 81434 79994
rect 81434 79942 81436 79994
rect 81380 79940 81436 79942
rect 81484 79994 81540 79996
rect 81484 79942 81486 79994
rect 81486 79942 81538 79994
rect 81538 79942 81540 79994
rect 81484 79940 81540 79942
rect 81276 78426 81332 78428
rect 81276 78374 81278 78426
rect 81278 78374 81330 78426
rect 81330 78374 81332 78426
rect 81276 78372 81332 78374
rect 81380 78426 81436 78428
rect 81380 78374 81382 78426
rect 81382 78374 81434 78426
rect 81434 78374 81436 78426
rect 81380 78372 81436 78374
rect 81484 78426 81540 78428
rect 81484 78374 81486 78426
rect 81486 78374 81538 78426
rect 81538 78374 81540 78426
rect 81484 78372 81540 78374
rect 81276 76858 81332 76860
rect 81276 76806 81278 76858
rect 81278 76806 81330 76858
rect 81330 76806 81332 76858
rect 81276 76804 81332 76806
rect 81380 76858 81436 76860
rect 81380 76806 81382 76858
rect 81382 76806 81434 76858
rect 81434 76806 81436 76858
rect 81380 76804 81436 76806
rect 81484 76858 81540 76860
rect 81484 76806 81486 76858
rect 81486 76806 81538 76858
rect 81538 76806 81540 76858
rect 81484 76804 81540 76806
rect 81276 75290 81332 75292
rect 81276 75238 81278 75290
rect 81278 75238 81330 75290
rect 81330 75238 81332 75290
rect 81276 75236 81332 75238
rect 81380 75290 81436 75292
rect 81380 75238 81382 75290
rect 81382 75238 81434 75290
rect 81434 75238 81436 75290
rect 81380 75236 81436 75238
rect 81484 75290 81540 75292
rect 81484 75238 81486 75290
rect 81486 75238 81538 75290
rect 81538 75238 81540 75290
rect 81484 75236 81540 75238
rect 81276 73722 81332 73724
rect 81276 73670 81278 73722
rect 81278 73670 81330 73722
rect 81330 73670 81332 73722
rect 81276 73668 81332 73670
rect 81380 73722 81436 73724
rect 81380 73670 81382 73722
rect 81382 73670 81434 73722
rect 81434 73670 81436 73722
rect 81380 73668 81436 73670
rect 81484 73722 81540 73724
rect 81484 73670 81486 73722
rect 81486 73670 81538 73722
rect 81538 73670 81540 73722
rect 81484 73668 81540 73670
rect 81276 72154 81332 72156
rect 81276 72102 81278 72154
rect 81278 72102 81330 72154
rect 81330 72102 81332 72154
rect 81276 72100 81332 72102
rect 81380 72154 81436 72156
rect 81380 72102 81382 72154
rect 81382 72102 81434 72154
rect 81434 72102 81436 72154
rect 81380 72100 81436 72102
rect 81484 72154 81540 72156
rect 81484 72102 81486 72154
rect 81486 72102 81538 72154
rect 81538 72102 81540 72154
rect 81484 72100 81540 72102
rect 81276 70586 81332 70588
rect 81276 70534 81278 70586
rect 81278 70534 81330 70586
rect 81330 70534 81332 70586
rect 81276 70532 81332 70534
rect 81380 70586 81436 70588
rect 81380 70534 81382 70586
rect 81382 70534 81434 70586
rect 81434 70534 81436 70586
rect 81380 70532 81436 70534
rect 81484 70586 81540 70588
rect 81484 70534 81486 70586
rect 81486 70534 81538 70586
rect 81538 70534 81540 70586
rect 81484 70532 81540 70534
rect 81276 69018 81332 69020
rect 81276 68966 81278 69018
rect 81278 68966 81330 69018
rect 81330 68966 81332 69018
rect 81276 68964 81332 68966
rect 81380 69018 81436 69020
rect 81380 68966 81382 69018
rect 81382 68966 81434 69018
rect 81434 68966 81436 69018
rect 81380 68964 81436 68966
rect 81484 69018 81540 69020
rect 81484 68966 81486 69018
rect 81486 68966 81538 69018
rect 81538 68966 81540 69018
rect 81484 68964 81540 68966
rect 81276 67450 81332 67452
rect 81276 67398 81278 67450
rect 81278 67398 81330 67450
rect 81330 67398 81332 67450
rect 81276 67396 81332 67398
rect 81380 67450 81436 67452
rect 81380 67398 81382 67450
rect 81382 67398 81434 67450
rect 81434 67398 81436 67450
rect 81380 67396 81436 67398
rect 81484 67450 81540 67452
rect 81484 67398 81486 67450
rect 81486 67398 81538 67450
rect 81538 67398 81540 67450
rect 81484 67396 81540 67398
rect 81276 65882 81332 65884
rect 81276 65830 81278 65882
rect 81278 65830 81330 65882
rect 81330 65830 81332 65882
rect 81276 65828 81332 65830
rect 81380 65882 81436 65884
rect 81380 65830 81382 65882
rect 81382 65830 81434 65882
rect 81434 65830 81436 65882
rect 81380 65828 81436 65830
rect 81484 65882 81540 65884
rect 81484 65830 81486 65882
rect 81486 65830 81538 65882
rect 81538 65830 81540 65882
rect 81484 65828 81540 65830
rect 81276 64314 81332 64316
rect 81276 64262 81278 64314
rect 81278 64262 81330 64314
rect 81330 64262 81332 64314
rect 81276 64260 81332 64262
rect 81380 64314 81436 64316
rect 81380 64262 81382 64314
rect 81382 64262 81434 64314
rect 81434 64262 81436 64314
rect 81380 64260 81436 64262
rect 81484 64314 81540 64316
rect 81484 64262 81486 64314
rect 81486 64262 81538 64314
rect 81538 64262 81540 64314
rect 81484 64260 81540 64262
rect 81276 62746 81332 62748
rect 81276 62694 81278 62746
rect 81278 62694 81330 62746
rect 81330 62694 81332 62746
rect 81276 62692 81332 62694
rect 81380 62746 81436 62748
rect 81380 62694 81382 62746
rect 81382 62694 81434 62746
rect 81434 62694 81436 62746
rect 81380 62692 81436 62694
rect 81484 62746 81540 62748
rect 81484 62694 81486 62746
rect 81486 62694 81538 62746
rect 81538 62694 81540 62746
rect 81484 62692 81540 62694
rect 81276 61178 81332 61180
rect 81276 61126 81278 61178
rect 81278 61126 81330 61178
rect 81330 61126 81332 61178
rect 81276 61124 81332 61126
rect 81380 61178 81436 61180
rect 81380 61126 81382 61178
rect 81382 61126 81434 61178
rect 81434 61126 81436 61178
rect 81380 61124 81436 61126
rect 81484 61178 81540 61180
rect 81484 61126 81486 61178
rect 81486 61126 81538 61178
rect 81538 61126 81540 61178
rect 81484 61124 81540 61126
rect 81276 59610 81332 59612
rect 81276 59558 81278 59610
rect 81278 59558 81330 59610
rect 81330 59558 81332 59610
rect 81276 59556 81332 59558
rect 81380 59610 81436 59612
rect 81380 59558 81382 59610
rect 81382 59558 81434 59610
rect 81434 59558 81436 59610
rect 81380 59556 81436 59558
rect 81484 59610 81540 59612
rect 81484 59558 81486 59610
rect 81486 59558 81538 59610
rect 81538 59558 81540 59610
rect 81484 59556 81540 59558
rect 81276 58042 81332 58044
rect 81276 57990 81278 58042
rect 81278 57990 81330 58042
rect 81330 57990 81332 58042
rect 81276 57988 81332 57990
rect 81380 58042 81436 58044
rect 81380 57990 81382 58042
rect 81382 57990 81434 58042
rect 81434 57990 81436 58042
rect 81380 57988 81436 57990
rect 81484 58042 81540 58044
rect 81484 57990 81486 58042
rect 81486 57990 81538 58042
rect 81538 57990 81540 58042
rect 81484 57988 81540 57990
rect 81276 56474 81332 56476
rect 81276 56422 81278 56474
rect 81278 56422 81330 56474
rect 81330 56422 81332 56474
rect 81276 56420 81332 56422
rect 81380 56474 81436 56476
rect 81380 56422 81382 56474
rect 81382 56422 81434 56474
rect 81434 56422 81436 56474
rect 81380 56420 81436 56422
rect 81484 56474 81540 56476
rect 81484 56422 81486 56474
rect 81486 56422 81538 56474
rect 81538 56422 81540 56474
rect 81484 56420 81540 56422
rect 81276 54906 81332 54908
rect 81276 54854 81278 54906
rect 81278 54854 81330 54906
rect 81330 54854 81332 54906
rect 81276 54852 81332 54854
rect 81380 54906 81436 54908
rect 81380 54854 81382 54906
rect 81382 54854 81434 54906
rect 81434 54854 81436 54906
rect 81380 54852 81436 54854
rect 81484 54906 81540 54908
rect 81484 54854 81486 54906
rect 81486 54854 81538 54906
rect 81538 54854 81540 54906
rect 81484 54852 81540 54854
rect 81276 53338 81332 53340
rect 81276 53286 81278 53338
rect 81278 53286 81330 53338
rect 81330 53286 81332 53338
rect 81276 53284 81332 53286
rect 81380 53338 81436 53340
rect 81380 53286 81382 53338
rect 81382 53286 81434 53338
rect 81434 53286 81436 53338
rect 81380 53284 81436 53286
rect 81484 53338 81540 53340
rect 81484 53286 81486 53338
rect 81486 53286 81538 53338
rect 81538 53286 81540 53338
rect 81484 53284 81540 53286
rect 81276 51770 81332 51772
rect 81276 51718 81278 51770
rect 81278 51718 81330 51770
rect 81330 51718 81332 51770
rect 81276 51716 81332 51718
rect 81380 51770 81436 51772
rect 81380 51718 81382 51770
rect 81382 51718 81434 51770
rect 81434 51718 81436 51770
rect 81380 51716 81436 51718
rect 81484 51770 81540 51772
rect 81484 51718 81486 51770
rect 81486 51718 81538 51770
rect 81538 51718 81540 51770
rect 81484 51716 81540 51718
rect 81276 50202 81332 50204
rect 81276 50150 81278 50202
rect 81278 50150 81330 50202
rect 81330 50150 81332 50202
rect 81276 50148 81332 50150
rect 81380 50202 81436 50204
rect 81380 50150 81382 50202
rect 81382 50150 81434 50202
rect 81434 50150 81436 50202
rect 81380 50148 81436 50150
rect 81484 50202 81540 50204
rect 81484 50150 81486 50202
rect 81486 50150 81538 50202
rect 81538 50150 81540 50202
rect 81484 50148 81540 50150
rect 81276 48634 81332 48636
rect 81276 48582 81278 48634
rect 81278 48582 81330 48634
rect 81330 48582 81332 48634
rect 81276 48580 81332 48582
rect 81380 48634 81436 48636
rect 81380 48582 81382 48634
rect 81382 48582 81434 48634
rect 81434 48582 81436 48634
rect 81380 48580 81436 48582
rect 81484 48634 81540 48636
rect 81484 48582 81486 48634
rect 81486 48582 81538 48634
rect 81538 48582 81540 48634
rect 81484 48580 81540 48582
rect 81276 47066 81332 47068
rect 81276 47014 81278 47066
rect 81278 47014 81330 47066
rect 81330 47014 81332 47066
rect 81276 47012 81332 47014
rect 81380 47066 81436 47068
rect 81380 47014 81382 47066
rect 81382 47014 81434 47066
rect 81434 47014 81436 47066
rect 81380 47012 81436 47014
rect 81484 47066 81540 47068
rect 81484 47014 81486 47066
rect 81486 47014 81538 47066
rect 81538 47014 81540 47066
rect 81484 47012 81540 47014
rect 81276 45498 81332 45500
rect 81276 45446 81278 45498
rect 81278 45446 81330 45498
rect 81330 45446 81332 45498
rect 81276 45444 81332 45446
rect 81380 45498 81436 45500
rect 81380 45446 81382 45498
rect 81382 45446 81434 45498
rect 81434 45446 81436 45498
rect 81380 45444 81436 45446
rect 81484 45498 81540 45500
rect 81484 45446 81486 45498
rect 81486 45446 81538 45498
rect 81538 45446 81540 45498
rect 81484 45444 81540 45446
rect 81276 43930 81332 43932
rect 81276 43878 81278 43930
rect 81278 43878 81330 43930
rect 81330 43878 81332 43930
rect 81276 43876 81332 43878
rect 81380 43930 81436 43932
rect 81380 43878 81382 43930
rect 81382 43878 81434 43930
rect 81434 43878 81436 43930
rect 81380 43876 81436 43878
rect 81484 43930 81540 43932
rect 81484 43878 81486 43930
rect 81486 43878 81538 43930
rect 81538 43878 81540 43930
rect 81484 43876 81540 43878
rect 81276 42362 81332 42364
rect 81276 42310 81278 42362
rect 81278 42310 81330 42362
rect 81330 42310 81332 42362
rect 81276 42308 81332 42310
rect 81380 42362 81436 42364
rect 81380 42310 81382 42362
rect 81382 42310 81434 42362
rect 81434 42310 81436 42362
rect 81380 42308 81436 42310
rect 81484 42362 81540 42364
rect 81484 42310 81486 42362
rect 81486 42310 81538 42362
rect 81538 42310 81540 42362
rect 81484 42308 81540 42310
rect 81276 40794 81332 40796
rect 81276 40742 81278 40794
rect 81278 40742 81330 40794
rect 81330 40742 81332 40794
rect 81276 40740 81332 40742
rect 81380 40794 81436 40796
rect 81380 40742 81382 40794
rect 81382 40742 81434 40794
rect 81434 40742 81436 40794
rect 81380 40740 81436 40742
rect 81484 40794 81540 40796
rect 81484 40742 81486 40794
rect 81486 40742 81538 40794
rect 81538 40742 81540 40794
rect 81484 40740 81540 40742
rect 81276 39226 81332 39228
rect 81276 39174 81278 39226
rect 81278 39174 81330 39226
rect 81330 39174 81332 39226
rect 81276 39172 81332 39174
rect 81380 39226 81436 39228
rect 81380 39174 81382 39226
rect 81382 39174 81434 39226
rect 81434 39174 81436 39226
rect 81380 39172 81436 39174
rect 81484 39226 81540 39228
rect 81484 39174 81486 39226
rect 81486 39174 81538 39226
rect 81538 39174 81540 39226
rect 81484 39172 81540 39174
rect 81276 37658 81332 37660
rect 81276 37606 81278 37658
rect 81278 37606 81330 37658
rect 81330 37606 81332 37658
rect 81276 37604 81332 37606
rect 81380 37658 81436 37660
rect 81380 37606 81382 37658
rect 81382 37606 81434 37658
rect 81434 37606 81436 37658
rect 81380 37604 81436 37606
rect 81484 37658 81540 37660
rect 81484 37606 81486 37658
rect 81486 37606 81538 37658
rect 81538 37606 81540 37658
rect 81484 37604 81540 37606
rect 81276 36090 81332 36092
rect 81276 36038 81278 36090
rect 81278 36038 81330 36090
rect 81330 36038 81332 36090
rect 81276 36036 81332 36038
rect 81380 36090 81436 36092
rect 81380 36038 81382 36090
rect 81382 36038 81434 36090
rect 81434 36038 81436 36090
rect 81380 36036 81436 36038
rect 81484 36090 81540 36092
rect 81484 36038 81486 36090
rect 81486 36038 81538 36090
rect 81538 36038 81540 36090
rect 81484 36036 81540 36038
rect 81276 34522 81332 34524
rect 81276 34470 81278 34522
rect 81278 34470 81330 34522
rect 81330 34470 81332 34522
rect 81276 34468 81332 34470
rect 81380 34522 81436 34524
rect 81380 34470 81382 34522
rect 81382 34470 81434 34522
rect 81434 34470 81436 34522
rect 81380 34468 81436 34470
rect 81484 34522 81540 34524
rect 81484 34470 81486 34522
rect 81486 34470 81538 34522
rect 81538 34470 81540 34522
rect 81484 34468 81540 34470
rect 81276 32954 81332 32956
rect 81276 32902 81278 32954
rect 81278 32902 81330 32954
rect 81330 32902 81332 32954
rect 81276 32900 81332 32902
rect 81380 32954 81436 32956
rect 81380 32902 81382 32954
rect 81382 32902 81434 32954
rect 81434 32902 81436 32954
rect 81380 32900 81436 32902
rect 81484 32954 81540 32956
rect 81484 32902 81486 32954
rect 81486 32902 81538 32954
rect 81538 32902 81540 32954
rect 81484 32900 81540 32902
rect 81276 31386 81332 31388
rect 81276 31334 81278 31386
rect 81278 31334 81330 31386
rect 81330 31334 81332 31386
rect 81276 31332 81332 31334
rect 81380 31386 81436 31388
rect 81380 31334 81382 31386
rect 81382 31334 81434 31386
rect 81434 31334 81436 31386
rect 81380 31332 81436 31334
rect 81484 31386 81540 31388
rect 81484 31334 81486 31386
rect 81486 31334 81538 31386
rect 81538 31334 81540 31386
rect 81484 31332 81540 31334
rect 81276 29818 81332 29820
rect 81276 29766 81278 29818
rect 81278 29766 81330 29818
rect 81330 29766 81332 29818
rect 81276 29764 81332 29766
rect 81380 29818 81436 29820
rect 81380 29766 81382 29818
rect 81382 29766 81434 29818
rect 81434 29766 81436 29818
rect 81380 29764 81436 29766
rect 81484 29818 81540 29820
rect 81484 29766 81486 29818
rect 81486 29766 81538 29818
rect 81538 29766 81540 29818
rect 81484 29764 81540 29766
rect 81276 28250 81332 28252
rect 81276 28198 81278 28250
rect 81278 28198 81330 28250
rect 81330 28198 81332 28250
rect 81276 28196 81332 28198
rect 81380 28250 81436 28252
rect 81380 28198 81382 28250
rect 81382 28198 81434 28250
rect 81434 28198 81436 28250
rect 81380 28196 81436 28198
rect 81484 28250 81540 28252
rect 81484 28198 81486 28250
rect 81486 28198 81538 28250
rect 81538 28198 81540 28250
rect 81484 28196 81540 28198
rect 81276 26682 81332 26684
rect 81276 26630 81278 26682
rect 81278 26630 81330 26682
rect 81330 26630 81332 26682
rect 81276 26628 81332 26630
rect 81380 26682 81436 26684
rect 81380 26630 81382 26682
rect 81382 26630 81434 26682
rect 81434 26630 81436 26682
rect 81380 26628 81436 26630
rect 81484 26682 81540 26684
rect 81484 26630 81486 26682
rect 81486 26630 81538 26682
rect 81538 26630 81540 26682
rect 81484 26628 81540 26630
rect 96636 116842 96692 116844
rect 96636 116790 96638 116842
rect 96638 116790 96690 116842
rect 96690 116790 96692 116842
rect 96636 116788 96692 116790
rect 96740 116842 96796 116844
rect 96740 116790 96742 116842
rect 96742 116790 96794 116842
rect 96794 116790 96796 116842
rect 96740 116788 96796 116790
rect 96844 116842 96900 116844
rect 96844 116790 96846 116842
rect 96846 116790 96898 116842
rect 96898 116790 96900 116842
rect 96844 116788 96900 116790
rect 97020 116508 97076 116564
rect 97916 116562 97972 116564
rect 97916 116510 97918 116562
rect 97918 116510 97970 116562
rect 97970 116510 97972 116562
rect 97916 116508 97972 116510
rect 101724 116620 101780 116676
rect 102508 116620 102564 116676
rect 98588 116508 98644 116564
rect 100044 116562 100100 116564
rect 100044 116510 100046 116562
rect 100046 116510 100098 116562
rect 100098 116510 100100 116562
rect 100044 116508 100100 116510
rect 103292 116508 103348 116564
rect 104188 116562 104244 116564
rect 104188 116510 104190 116562
rect 104190 116510 104242 116562
rect 104242 116510 104244 116562
rect 104188 116508 104244 116510
rect 106428 116508 106484 116564
rect 93884 115724 93940 115780
rect 94444 115778 94500 115780
rect 94444 115726 94446 115778
rect 94446 115726 94498 115778
rect 94498 115726 94500 115778
rect 94444 115724 94500 115726
rect 91420 115612 91476 115668
rect 91980 115666 92036 115668
rect 91980 115614 91982 115666
rect 91982 115614 92034 115666
rect 92034 115614 92036 115666
rect 91980 115612 92036 115614
rect 96460 115666 96516 115668
rect 96460 115614 96462 115666
rect 96462 115614 96514 115666
rect 96514 115614 96516 115666
rect 96460 115612 96516 115614
rect 97580 115666 97636 115668
rect 97580 115614 97582 115666
rect 97582 115614 97634 115666
rect 97634 115614 97636 115666
rect 97580 115612 97636 115614
rect 100828 115666 100884 115668
rect 100828 115614 100830 115666
rect 100830 115614 100882 115666
rect 100882 115614 100884 115666
rect 100828 115612 100884 115614
rect 95340 115500 95396 115556
rect 95900 115554 95956 115556
rect 95900 115502 95902 115554
rect 95902 115502 95954 115554
rect 95954 115502 95956 115554
rect 95900 115500 95956 115502
rect 97468 115500 97524 115556
rect 96636 115274 96692 115276
rect 96636 115222 96638 115274
rect 96638 115222 96690 115274
rect 96690 115222 96692 115274
rect 96636 115220 96692 115222
rect 96740 115274 96796 115276
rect 96740 115222 96742 115274
rect 96742 115222 96794 115274
rect 96794 115222 96796 115274
rect 96740 115220 96796 115222
rect 96844 115274 96900 115276
rect 96844 115222 96846 115274
rect 96846 115222 96898 115274
rect 96898 115222 96900 115274
rect 96844 115220 96900 115222
rect 91420 114828 91476 114884
rect 96636 113706 96692 113708
rect 96636 113654 96638 113706
rect 96638 113654 96690 113706
rect 96690 113654 96692 113706
rect 96636 113652 96692 113654
rect 96740 113706 96796 113708
rect 96740 113654 96742 113706
rect 96742 113654 96794 113706
rect 96794 113654 96796 113706
rect 96740 113652 96796 113654
rect 96844 113706 96900 113708
rect 96844 113654 96846 113706
rect 96846 113654 96898 113706
rect 96898 113654 96900 113706
rect 96844 113652 96900 113654
rect 96636 112138 96692 112140
rect 96636 112086 96638 112138
rect 96638 112086 96690 112138
rect 96690 112086 96692 112138
rect 96636 112084 96692 112086
rect 96740 112138 96796 112140
rect 96740 112086 96742 112138
rect 96742 112086 96794 112138
rect 96794 112086 96796 112138
rect 96740 112084 96796 112086
rect 96844 112138 96900 112140
rect 96844 112086 96846 112138
rect 96846 112086 96898 112138
rect 96898 112086 96900 112138
rect 96844 112084 96900 112086
rect 96636 110570 96692 110572
rect 96636 110518 96638 110570
rect 96638 110518 96690 110570
rect 96690 110518 96692 110570
rect 96636 110516 96692 110518
rect 96740 110570 96796 110572
rect 96740 110518 96742 110570
rect 96742 110518 96794 110570
rect 96794 110518 96796 110570
rect 96740 110516 96796 110518
rect 96844 110570 96900 110572
rect 96844 110518 96846 110570
rect 96846 110518 96898 110570
rect 96898 110518 96900 110570
rect 96844 110516 96900 110518
rect 96636 109002 96692 109004
rect 96636 108950 96638 109002
rect 96638 108950 96690 109002
rect 96690 108950 96692 109002
rect 96636 108948 96692 108950
rect 96740 109002 96796 109004
rect 96740 108950 96742 109002
rect 96742 108950 96794 109002
rect 96794 108950 96796 109002
rect 96740 108948 96796 108950
rect 96844 109002 96900 109004
rect 96844 108950 96846 109002
rect 96846 108950 96898 109002
rect 96898 108950 96900 109002
rect 96844 108948 96900 108950
rect 96636 107434 96692 107436
rect 96636 107382 96638 107434
rect 96638 107382 96690 107434
rect 96690 107382 96692 107434
rect 96636 107380 96692 107382
rect 96740 107434 96796 107436
rect 96740 107382 96742 107434
rect 96742 107382 96794 107434
rect 96794 107382 96796 107434
rect 96740 107380 96796 107382
rect 96844 107434 96900 107436
rect 96844 107382 96846 107434
rect 96846 107382 96898 107434
rect 96898 107382 96900 107434
rect 96844 107380 96900 107382
rect 96636 105866 96692 105868
rect 96636 105814 96638 105866
rect 96638 105814 96690 105866
rect 96690 105814 96692 105866
rect 96636 105812 96692 105814
rect 96740 105866 96796 105868
rect 96740 105814 96742 105866
rect 96742 105814 96794 105866
rect 96794 105814 96796 105866
rect 96740 105812 96796 105814
rect 96844 105866 96900 105868
rect 96844 105814 96846 105866
rect 96846 105814 96898 105866
rect 96898 105814 96900 105866
rect 96844 105812 96900 105814
rect 96636 104298 96692 104300
rect 96636 104246 96638 104298
rect 96638 104246 96690 104298
rect 96690 104246 96692 104298
rect 96636 104244 96692 104246
rect 96740 104298 96796 104300
rect 96740 104246 96742 104298
rect 96742 104246 96794 104298
rect 96794 104246 96796 104298
rect 96740 104244 96796 104246
rect 96844 104298 96900 104300
rect 96844 104246 96846 104298
rect 96846 104246 96898 104298
rect 96898 104246 96900 104298
rect 96844 104244 96900 104246
rect 96636 102730 96692 102732
rect 96636 102678 96638 102730
rect 96638 102678 96690 102730
rect 96690 102678 96692 102730
rect 96636 102676 96692 102678
rect 96740 102730 96796 102732
rect 96740 102678 96742 102730
rect 96742 102678 96794 102730
rect 96794 102678 96796 102730
rect 96740 102676 96796 102678
rect 96844 102730 96900 102732
rect 96844 102678 96846 102730
rect 96846 102678 96898 102730
rect 96898 102678 96900 102730
rect 96844 102676 96900 102678
rect 96636 101162 96692 101164
rect 96636 101110 96638 101162
rect 96638 101110 96690 101162
rect 96690 101110 96692 101162
rect 96636 101108 96692 101110
rect 96740 101162 96796 101164
rect 96740 101110 96742 101162
rect 96742 101110 96794 101162
rect 96794 101110 96796 101162
rect 96740 101108 96796 101110
rect 96844 101162 96900 101164
rect 96844 101110 96846 101162
rect 96846 101110 96898 101162
rect 96898 101110 96900 101162
rect 96844 101108 96900 101110
rect 96636 99594 96692 99596
rect 96636 99542 96638 99594
rect 96638 99542 96690 99594
rect 96690 99542 96692 99594
rect 96636 99540 96692 99542
rect 96740 99594 96796 99596
rect 96740 99542 96742 99594
rect 96742 99542 96794 99594
rect 96794 99542 96796 99594
rect 96740 99540 96796 99542
rect 96844 99594 96900 99596
rect 96844 99542 96846 99594
rect 96846 99542 96898 99594
rect 96898 99542 96900 99594
rect 96844 99540 96900 99542
rect 96636 98026 96692 98028
rect 96636 97974 96638 98026
rect 96638 97974 96690 98026
rect 96690 97974 96692 98026
rect 96636 97972 96692 97974
rect 96740 98026 96796 98028
rect 96740 97974 96742 98026
rect 96742 97974 96794 98026
rect 96794 97974 96796 98026
rect 96740 97972 96796 97974
rect 96844 98026 96900 98028
rect 96844 97974 96846 98026
rect 96846 97974 96898 98026
rect 96898 97974 96900 98026
rect 96844 97972 96900 97974
rect 96636 96458 96692 96460
rect 96636 96406 96638 96458
rect 96638 96406 96690 96458
rect 96690 96406 96692 96458
rect 96636 96404 96692 96406
rect 96740 96458 96796 96460
rect 96740 96406 96742 96458
rect 96742 96406 96794 96458
rect 96794 96406 96796 96458
rect 96740 96404 96796 96406
rect 96844 96458 96900 96460
rect 96844 96406 96846 96458
rect 96846 96406 96898 96458
rect 96898 96406 96900 96458
rect 96844 96404 96900 96406
rect 96636 94890 96692 94892
rect 96636 94838 96638 94890
rect 96638 94838 96690 94890
rect 96690 94838 96692 94890
rect 96636 94836 96692 94838
rect 96740 94890 96796 94892
rect 96740 94838 96742 94890
rect 96742 94838 96794 94890
rect 96794 94838 96796 94890
rect 96740 94836 96796 94838
rect 96844 94890 96900 94892
rect 96844 94838 96846 94890
rect 96846 94838 96898 94890
rect 96898 94838 96900 94890
rect 96844 94836 96900 94838
rect 96636 93322 96692 93324
rect 96636 93270 96638 93322
rect 96638 93270 96690 93322
rect 96690 93270 96692 93322
rect 96636 93268 96692 93270
rect 96740 93322 96796 93324
rect 96740 93270 96742 93322
rect 96742 93270 96794 93322
rect 96794 93270 96796 93322
rect 96740 93268 96796 93270
rect 96844 93322 96900 93324
rect 96844 93270 96846 93322
rect 96846 93270 96898 93322
rect 96898 93270 96900 93322
rect 96844 93268 96900 93270
rect 96636 91754 96692 91756
rect 96636 91702 96638 91754
rect 96638 91702 96690 91754
rect 96690 91702 96692 91754
rect 96636 91700 96692 91702
rect 96740 91754 96796 91756
rect 96740 91702 96742 91754
rect 96742 91702 96794 91754
rect 96794 91702 96796 91754
rect 96740 91700 96796 91702
rect 96844 91754 96900 91756
rect 96844 91702 96846 91754
rect 96846 91702 96898 91754
rect 96898 91702 96900 91754
rect 96844 91700 96900 91702
rect 96636 90186 96692 90188
rect 96636 90134 96638 90186
rect 96638 90134 96690 90186
rect 96690 90134 96692 90186
rect 96636 90132 96692 90134
rect 96740 90186 96796 90188
rect 96740 90134 96742 90186
rect 96742 90134 96794 90186
rect 96794 90134 96796 90186
rect 96740 90132 96796 90134
rect 96844 90186 96900 90188
rect 96844 90134 96846 90186
rect 96846 90134 96898 90186
rect 96898 90134 96900 90186
rect 96844 90132 96900 90134
rect 96636 88618 96692 88620
rect 96636 88566 96638 88618
rect 96638 88566 96690 88618
rect 96690 88566 96692 88618
rect 96636 88564 96692 88566
rect 96740 88618 96796 88620
rect 96740 88566 96742 88618
rect 96742 88566 96794 88618
rect 96794 88566 96796 88618
rect 96740 88564 96796 88566
rect 96844 88618 96900 88620
rect 96844 88566 96846 88618
rect 96846 88566 96898 88618
rect 96898 88566 96900 88618
rect 96844 88564 96900 88566
rect 96636 87050 96692 87052
rect 96636 86998 96638 87050
rect 96638 86998 96690 87050
rect 96690 86998 96692 87050
rect 96636 86996 96692 86998
rect 96740 87050 96796 87052
rect 96740 86998 96742 87050
rect 96742 86998 96794 87050
rect 96794 86998 96796 87050
rect 96740 86996 96796 86998
rect 96844 87050 96900 87052
rect 96844 86998 96846 87050
rect 96846 86998 96898 87050
rect 96898 86998 96900 87050
rect 96844 86996 96900 86998
rect 96636 85482 96692 85484
rect 96636 85430 96638 85482
rect 96638 85430 96690 85482
rect 96690 85430 96692 85482
rect 96636 85428 96692 85430
rect 96740 85482 96796 85484
rect 96740 85430 96742 85482
rect 96742 85430 96794 85482
rect 96794 85430 96796 85482
rect 96740 85428 96796 85430
rect 96844 85482 96900 85484
rect 96844 85430 96846 85482
rect 96846 85430 96898 85482
rect 96898 85430 96900 85482
rect 96844 85428 96900 85430
rect 96636 83914 96692 83916
rect 96636 83862 96638 83914
rect 96638 83862 96690 83914
rect 96690 83862 96692 83914
rect 96636 83860 96692 83862
rect 96740 83914 96796 83916
rect 96740 83862 96742 83914
rect 96742 83862 96794 83914
rect 96794 83862 96796 83914
rect 96740 83860 96796 83862
rect 96844 83914 96900 83916
rect 96844 83862 96846 83914
rect 96846 83862 96898 83914
rect 96898 83862 96900 83914
rect 96844 83860 96900 83862
rect 96636 82346 96692 82348
rect 96636 82294 96638 82346
rect 96638 82294 96690 82346
rect 96690 82294 96692 82346
rect 96636 82292 96692 82294
rect 96740 82346 96796 82348
rect 96740 82294 96742 82346
rect 96742 82294 96794 82346
rect 96794 82294 96796 82346
rect 96740 82292 96796 82294
rect 96844 82346 96900 82348
rect 96844 82294 96846 82346
rect 96846 82294 96898 82346
rect 96898 82294 96900 82346
rect 96844 82292 96900 82294
rect 96636 80778 96692 80780
rect 96636 80726 96638 80778
rect 96638 80726 96690 80778
rect 96690 80726 96692 80778
rect 96636 80724 96692 80726
rect 96740 80778 96796 80780
rect 96740 80726 96742 80778
rect 96742 80726 96794 80778
rect 96794 80726 96796 80778
rect 96740 80724 96796 80726
rect 96844 80778 96900 80780
rect 96844 80726 96846 80778
rect 96846 80726 96898 80778
rect 96898 80726 96900 80778
rect 96844 80724 96900 80726
rect 96636 79210 96692 79212
rect 96636 79158 96638 79210
rect 96638 79158 96690 79210
rect 96690 79158 96692 79210
rect 96636 79156 96692 79158
rect 96740 79210 96796 79212
rect 96740 79158 96742 79210
rect 96742 79158 96794 79210
rect 96794 79158 96796 79210
rect 96740 79156 96796 79158
rect 96844 79210 96900 79212
rect 96844 79158 96846 79210
rect 96846 79158 96898 79210
rect 96898 79158 96900 79210
rect 96844 79156 96900 79158
rect 96636 77642 96692 77644
rect 96636 77590 96638 77642
rect 96638 77590 96690 77642
rect 96690 77590 96692 77642
rect 96636 77588 96692 77590
rect 96740 77642 96796 77644
rect 96740 77590 96742 77642
rect 96742 77590 96794 77642
rect 96794 77590 96796 77642
rect 96740 77588 96796 77590
rect 96844 77642 96900 77644
rect 96844 77590 96846 77642
rect 96846 77590 96898 77642
rect 96898 77590 96900 77642
rect 96844 77588 96900 77590
rect 96636 76074 96692 76076
rect 96636 76022 96638 76074
rect 96638 76022 96690 76074
rect 96690 76022 96692 76074
rect 96636 76020 96692 76022
rect 96740 76074 96796 76076
rect 96740 76022 96742 76074
rect 96742 76022 96794 76074
rect 96794 76022 96796 76074
rect 96740 76020 96796 76022
rect 96844 76074 96900 76076
rect 96844 76022 96846 76074
rect 96846 76022 96898 76074
rect 96898 76022 96900 76074
rect 96844 76020 96900 76022
rect 96636 74506 96692 74508
rect 96636 74454 96638 74506
rect 96638 74454 96690 74506
rect 96690 74454 96692 74506
rect 96636 74452 96692 74454
rect 96740 74506 96796 74508
rect 96740 74454 96742 74506
rect 96742 74454 96794 74506
rect 96794 74454 96796 74506
rect 96740 74452 96796 74454
rect 96844 74506 96900 74508
rect 96844 74454 96846 74506
rect 96846 74454 96898 74506
rect 96898 74454 96900 74506
rect 96844 74452 96900 74454
rect 96636 72938 96692 72940
rect 96636 72886 96638 72938
rect 96638 72886 96690 72938
rect 96690 72886 96692 72938
rect 96636 72884 96692 72886
rect 96740 72938 96796 72940
rect 96740 72886 96742 72938
rect 96742 72886 96794 72938
rect 96794 72886 96796 72938
rect 96740 72884 96796 72886
rect 96844 72938 96900 72940
rect 96844 72886 96846 72938
rect 96846 72886 96898 72938
rect 96898 72886 96900 72938
rect 96844 72884 96900 72886
rect 96636 71370 96692 71372
rect 96636 71318 96638 71370
rect 96638 71318 96690 71370
rect 96690 71318 96692 71370
rect 96636 71316 96692 71318
rect 96740 71370 96796 71372
rect 96740 71318 96742 71370
rect 96742 71318 96794 71370
rect 96794 71318 96796 71370
rect 96740 71316 96796 71318
rect 96844 71370 96900 71372
rect 96844 71318 96846 71370
rect 96846 71318 96898 71370
rect 96898 71318 96900 71370
rect 96844 71316 96900 71318
rect 96636 69802 96692 69804
rect 96636 69750 96638 69802
rect 96638 69750 96690 69802
rect 96690 69750 96692 69802
rect 96636 69748 96692 69750
rect 96740 69802 96796 69804
rect 96740 69750 96742 69802
rect 96742 69750 96794 69802
rect 96794 69750 96796 69802
rect 96740 69748 96796 69750
rect 96844 69802 96900 69804
rect 96844 69750 96846 69802
rect 96846 69750 96898 69802
rect 96898 69750 96900 69802
rect 96844 69748 96900 69750
rect 96636 68234 96692 68236
rect 96636 68182 96638 68234
rect 96638 68182 96690 68234
rect 96690 68182 96692 68234
rect 96636 68180 96692 68182
rect 96740 68234 96796 68236
rect 96740 68182 96742 68234
rect 96742 68182 96794 68234
rect 96794 68182 96796 68234
rect 96740 68180 96796 68182
rect 96844 68234 96900 68236
rect 96844 68182 96846 68234
rect 96846 68182 96898 68234
rect 96898 68182 96900 68234
rect 96844 68180 96900 68182
rect 96636 66666 96692 66668
rect 96636 66614 96638 66666
rect 96638 66614 96690 66666
rect 96690 66614 96692 66666
rect 96636 66612 96692 66614
rect 96740 66666 96796 66668
rect 96740 66614 96742 66666
rect 96742 66614 96794 66666
rect 96794 66614 96796 66666
rect 96740 66612 96796 66614
rect 96844 66666 96900 66668
rect 96844 66614 96846 66666
rect 96846 66614 96898 66666
rect 96898 66614 96900 66666
rect 96844 66612 96900 66614
rect 96636 65098 96692 65100
rect 96636 65046 96638 65098
rect 96638 65046 96690 65098
rect 96690 65046 96692 65098
rect 96636 65044 96692 65046
rect 96740 65098 96796 65100
rect 96740 65046 96742 65098
rect 96742 65046 96794 65098
rect 96794 65046 96796 65098
rect 96740 65044 96796 65046
rect 96844 65098 96900 65100
rect 96844 65046 96846 65098
rect 96846 65046 96898 65098
rect 96898 65046 96900 65098
rect 96844 65044 96900 65046
rect 96636 63530 96692 63532
rect 96636 63478 96638 63530
rect 96638 63478 96690 63530
rect 96690 63478 96692 63530
rect 96636 63476 96692 63478
rect 96740 63530 96796 63532
rect 96740 63478 96742 63530
rect 96742 63478 96794 63530
rect 96794 63478 96796 63530
rect 96740 63476 96796 63478
rect 96844 63530 96900 63532
rect 96844 63478 96846 63530
rect 96846 63478 96898 63530
rect 96898 63478 96900 63530
rect 96844 63476 96900 63478
rect 96636 61962 96692 61964
rect 96636 61910 96638 61962
rect 96638 61910 96690 61962
rect 96690 61910 96692 61962
rect 96636 61908 96692 61910
rect 96740 61962 96796 61964
rect 96740 61910 96742 61962
rect 96742 61910 96794 61962
rect 96794 61910 96796 61962
rect 96740 61908 96796 61910
rect 96844 61962 96900 61964
rect 96844 61910 96846 61962
rect 96846 61910 96898 61962
rect 96898 61910 96900 61962
rect 96844 61908 96900 61910
rect 96636 60394 96692 60396
rect 96636 60342 96638 60394
rect 96638 60342 96690 60394
rect 96690 60342 96692 60394
rect 96636 60340 96692 60342
rect 96740 60394 96796 60396
rect 96740 60342 96742 60394
rect 96742 60342 96794 60394
rect 96794 60342 96796 60394
rect 96740 60340 96796 60342
rect 96844 60394 96900 60396
rect 96844 60342 96846 60394
rect 96846 60342 96898 60394
rect 96898 60342 96900 60394
rect 96844 60340 96900 60342
rect 96636 58826 96692 58828
rect 96636 58774 96638 58826
rect 96638 58774 96690 58826
rect 96690 58774 96692 58826
rect 96636 58772 96692 58774
rect 96740 58826 96796 58828
rect 96740 58774 96742 58826
rect 96742 58774 96794 58826
rect 96794 58774 96796 58826
rect 96740 58772 96796 58774
rect 96844 58826 96900 58828
rect 96844 58774 96846 58826
rect 96846 58774 96898 58826
rect 96898 58774 96900 58826
rect 96844 58772 96900 58774
rect 96636 57258 96692 57260
rect 96636 57206 96638 57258
rect 96638 57206 96690 57258
rect 96690 57206 96692 57258
rect 96636 57204 96692 57206
rect 96740 57258 96796 57260
rect 96740 57206 96742 57258
rect 96742 57206 96794 57258
rect 96794 57206 96796 57258
rect 96740 57204 96796 57206
rect 96844 57258 96900 57260
rect 96844 57206 96846 57258
rect 96846 57206 96898 57258
rect 96898 57206 96900 57258
rect 96844 57204 96900 57206
rect 96636 55690 96692 55692
rect 96636 55638 96638 55690
rect 96638 55638 96690 55690
rect 96690 55638 96692 55690
rect 96636 55636 96692 55638
rect 96740 55690 96796 55692
rect 96740 55638 96742 55690
rect 96742 55638 96794 55690
rect 96794 55638 96796 55690
rect 96740 55636 96796 55638
rect 96844 55690 96900 55692
rect 96844 55638 96846 55690
rect 96846 55638 96898 55690
rect 96898 55638 96900 55690
rect 96844 55636 96900 55638
rect 96636 54122 96692 54124
rect 96636 54070 96638 54122
rect 96638 54070 96690 54122
rect 96690 54070 96692 54122
rect 96636 54068 96692 54070
rect 96740 54122 96796 54124
rect 96740 54070 96742 54122
rect 96742 54070 96794 54122
rect 96794 54070 96796 54122
rect 96740 54068 96796 54070
rect 96844 54122 96900 54124
rect 96844 54070 96846 54122
rect 96846 54070 96898 54122
rect 96898 54070 96900 54122
rect 96844 54068 96900 54070
rect 96636 52554 96692 52556
rect 96636 52502 96638 52554
rect 96638 52502 96690 52554
rect 96690 52502 96692 52554
rect 96636 52500 96692 52502
rect 96740 52554 96796 52556
rect 96740 52502 96742 52554
rect 96742 52502 96794 52554
rect 96794 52502 96796 52554
rect 96740 52500 96796 52502
rect 96844 52554 96900 52556
rect 96844 52502 96846 52554
rect 96846 52502 96898 52554
rect 96898 52502 96900 52554
rect 96844 52500 96900 52502
rect 96636 50986 96692 50988
rect 96636 50934 96638 50986
rect 96638 50934 96690 50986
rect 96690 50934 96692 50986
rect 96636 50932 96692 50934
rect 96740 50986 96796 50988
rect 96740 50934 96742 50986
rect 96742 50934 96794 50986
rect 96794 50934 96796 50986
rect 96740 50932 96796 50934
rect 96844 50986 96900 50988
rect 96844 50934 96846 50986
rect 96846 50934 96898 50986
rect 96898 50934 96900 50986
rect 96844 50932 96900 50934
rect 96636 49418 96692 49420
rect 96636 49366 96638 49418
rect 96638 49366 96690 49418
rect 96690 49366 96692 49418
rect 96636 49364 96692 49366
rect 96740 49418 96796 49420
rect 96740 49366 96742 49418
rect 96742 49366 96794 49418
rect 96794 49366 96796 49418
rect 96740 49364 96796 49366
rect 96844 49418 96900 49420
rect 96844 49366 96846 49418
rect 96846 49366 96898 49418
rect 96898 49366 96900 49418
rect 96844 49364 96900 49366
rect 96636 47850 96692 47852
rect 96636 47798 96638 47850
rect 96638 47798 96690 47850
rect 96690 47798 96692 47850
rect 96636 47796 96692 47798
rect 96740 47850 96796 47852
rect 96740 47798 96742 47850
rect 96742 47798 96794 47850
rect 96794 47798 96796 47850
rect 96740 47796 96796 47798
rect 96844 47850 96900 47852
rect 96844 47798 96846 47850
rect 96846 47798 96898 47850
rect 96898 47798 96900 47850
rect 96844 47796 96900 47798
rect 96636 46282 96692 46284
rect 96636 46230 96638 46282
rect 96638 46230 96690 46282
rect 96690 46230 96692 46282
rect 96636 46228 96692 46230
rect 96740 46282 96796 46284
rect 96740 46230 96742 46282
rect 96742 46230 96794 46282
rect 96794 46230 96796 46282
rect 96740 46228 96796 46230
rect 96844 46282 96900 46284
rect 96844 46230 96846 46282
rect 96846 46230 96898 46282
rect 96898 46230 96900 46282
rect 96844 46228 96900 46230
rect 96636 44714 96692 44716
rect 96636 44662 96638 44714
rect 96638 44662 96690 44714
rect 96690 44662 96692 44714
rect 96636 44660 96692 44662
rect 96740 44714 96796 44716
rect 96740 44662 96742 44714
rect 96742 44662 96794 44714
rect 96794 44662 96796 44714
rect 96740 44660 96796 44662
rect 96844 44714 96900 44716
rect 96844 44662 96846 44714
rect 96846 44662 96898 44714
rect 96898 44662 96900 44714
rect 96844 44660 96900 44662
rect 96636 43146 96692 43148
rect 96636 43094 96638 43146
rect 96638 43094 96690 43146
rect 96690 43094 96692 43146
rect 96636 43092 96692 43094
rect 96740 43146 96796 43148
rect 96740 43094 96742 43146
rect 96742 43094 96794 43146
rect 96794 43094 96796 43146
rect 96740 43092 96796 43094
rect 96844 43146 96900 43148
rect 96844 43094 96846 43146
rect 96846 43094 96898 43146
rect 96898 43094 96900 43146
rect 96844 43092 96900 43094
rect 96636 41578 96692 41580
rect 96636 41526 96638 41578
rect 96638 41526 96690 41578
rect 96690 41526 96692 41578
rect 96636 41524 96692 41526
rect 96740 41578 96796 41580
rect 96740 41526 96742 41578
rect 96742 41526 96794 41578
rect 96794 41526 96796 41578
rect 96740 41524 96796 41526
rect 96844 41578 96900 41580
rect 96844 41526 96846 41578
rect 96846 41526 96898 41578
rect 96898 41526 96900 41578
rect 96844 41524 96900 41526
rect 96636 40010 96692 40012
rect 96636 39958 96638 40010
rect 96638 39958 96690 40010
rect 96690 39958 96692 40010
rect 96636 39956 96692 39958
rect 96740 40010 96796 40012
rect 96740 39958 96742 40010
rect 96742 39958 96794 40010
rect 96794 39958 96796 40010
rect 96740 39956 96796 39958
rect 96844 40010 96900 40012
rect 96844 39958 96846 40010
rect 96846 39958 96898 40010
rect 96898 39958 96900 40010
rect 96844 39956 96900 39958
rect 96636 38442 96692 38444
rect 96636 38390 96638 38442
rect 96638 38390 96690 38442
rect 96690 38390 96692 38442
rect 96636 38388 96692 38390
rect 96740 38442 96796 38444
rect 96740 38390 96742 38442
rect 96742 38390 96794 38442
rect 96794 38390 96796 38442
rect 96740 38388 96796 38390
rect 96844 38442 96900 38444
rect 96844 38390 96846 38442
rect 96846 38390 96898 38442
rect 96898 38390 96900 38442
rect 96844 38388 96900 38390
rect 96636 36874 96692 36876
rect 96636 36822 96638 36874
rect 96638 36822 96690 36874
rect 96690 36822 96692 36874
rect 96636 36820 96692 36822
rect 96740 36874 96796 36876
rect 96740 36822 96742 36874
rect 96742 36822 96794 36874
rect 96794 36822 96796 36874
rect 96740 36820 96796 36822
rect 96844 36874 96900 36876
rect 96844 36822 96846 36874
rect 96846 36822 96898 36874
rect 96898 36822 96900 36874
rect 96844 36820 96900 36822
rect 96636 35306 96692 35308
rect 96636 35254 96638 35306
rect 96638 35254 96690 35306
rect 96690 35254 96692 35306
rect 96636 35252 96692 35254
rect 96740 35306 96796 35308
rect 96740 35254 96742 35306
rect 96742 35254 96794 35306
rect 96794 35254 96796 35306
rect 96740 35252 96796 35254
rect 96844 35306 96900 35308
rect 96844 35254 96846 35306
rect 96846 35254 96898 35306
rect 96898 35254 96900 35306
rect 96844 35252 96900 35254
rect 96636 33738 96692 33740
rect 96636 33686 96638 33738
rect 96638 33686 96690 33738
rect 96690 33686 96692 33738
rect 96636 33684 96692 33686
rect 96740 33738 96796 33740
rect 96740 33686 96742 33738
rect 96742 33686 96794 33738
rect 96794 33686 96796 33738
rect 96740 33684 96796 33686
rect 96844 33738 96900 33740
rect 96844 33686 96846 33738
rect 96846 33686 96898 33738
rect 96898 33686 96900 33738
rect 96844 33684 96900 33686
rect 96636 32170 96692 32172
rect 96636 32118 96638 32170
rect 96638 32118 96690 32170
rect 96690 32118 96692 32170
rect 96636 32116 96692 32118
rect 96740 32170 96796 32172
rect 96740 32118 96742 32170
rect 96742 32118 96794 32170
rect 96794 32118 96796 32170
rect 96740 32116 96796 32118
rect 96844 32170 96900 32172
rect 96844 32118 96846 32170
rect 96846 32118 96898 32170
rect 96898 32118 96900 32170
rect 96844 32116 96900 32118
rect 96636 30602 96692 30604
rect 96636 30550 96638 30602
rect 96638 30550 96690 30602
rect 96690 30550 96692 30602
rect 96636 30548 96692 30550
rect 96740 30602 96796 30604
rect 96740 30550 96742 30602
rect 96742 30550 96794 30602
rect 96794 30550 96796 30602
rect 96740 30548 96796 30550
rect 96844 30602 96900 30604
rect 96844 30550 96846 30602
rect 96846 30550 96898 30602
rect 96898 30550 96900 30602
rect 96844 30548 96900 30550
rect 96636 29034 96692 29036
rect 96636 28982 96638 29034
rect 96638 28982 96690 29034
rect 96690 28982 96692 29034
rect 96636 28980 96692 28982
rect 96740 29034 96796 29036
rect 96740 28982 96742 29034
rect 96742 28982 96794 29034
rect 96794 28982 96796 29034
rect 96740 28980 96796 28982
rect 96844 29034 96900 29036
rect 96844 28982 96846 29034
rect 96846 28982 96898 29034
rect 96898 28982 96900 29034
rect 96844 28980 96900 28982
rect 96636 27466 96692 27468
rect 96636 27414 96638 27466
rect 96638 27414 96690 27466
rect 96690 27414 96692 27466
rect 96636 27412 96692 27414
rect 96740 27466 96796 27468
rect 96740 27414 96742 27466
rect 96742 27414 96794 27466
rect 96794 27414 96796 27466
rect 96740 27412 96796 27414
rect 96844 27466 96900 27468
rect 96844 27414 96846 27466
rect 96846 27414 96898 27466
rect 96898 27414 96900 27466
rect 96844 27412 96900 27414
rect 106316 116396 106372 116452
rect 104972 116172 105028 116228
rect 105420 116226 105476 116228
rect 105420 116174 105422 116226
rect 105422 116174 105474 116226
rect 105474 116174 105476 116226
rect 105420 116172 105476 116174
rect 106092 116172 106148 116228
rect 101388 115666 101444 115668
rect 101388 115614 101390 115666
rect 101390 115614 101442 115666
rect 101442 115614 101444 115666
rect 101388 115612 101444 115614
rect 105420 115666 105476 115668
rect 105420 115614 105422 115666
rect 105422 115614 105474 115666
rect 105474 115614 105476 115666
rect 105420 115612 105476 115614
rect 105980 115666 106036 115668
rect 105980 115614 105982 115666
rect 105982 115614 106034 115666
rect 106034 115614 106036 115666
rect 105980 115612 106036 115614
rect 97468 27244 97524 27300
rect 98364 27244 98420 27300
rect 96636 25898 96692 25900
rect 96636 25846 96638 25898
rect 96638 25846 96690 25898
rect 96690 25846 96692 25898
rect 96636 25844 96692 25846
rect 96740 25898 96796 25900
rect 96740 25846 96742 25898
rect 96742 25846 96794 25898
rect 96794 25846 96796 25898
rect 96740 25844 96796 25846
rect 96844 25898 96900 25900
rect 96844 25846 96846 25898
rect 96846 25846 96898 25898
rect 96898 25846 96900 25898
rect 96844 25844 96900 25846
rect 90860 25564 90916 25620
rect 91532 25564 91588 25620
rect 81276 25114 81332 25116
rect 81276 25062 81278 25114
rect 81278 25062 81330 25114
rect 81330 25062 81332 25114
rect 81276 25060 81332 25062
rect 81380 25114 81436 25116
rect 81380 25062 81382 25114
rect 81382 25062 81434 25114
rect 81434 25062 81436 25114
rect 81380 25060 81436 25062
rect 81484 25114 81540 25116
rect 81484 25062 81486 25114
rect 81486 25062 81538 25114
rect 81538 25062 81540 25114
rect 81484 25060 81540 25062
rect 81276 23546 81332 23548
rect 81276 23494 81278 23546
rect 81278 23494 81330 23546
rect 81330 23494 81332 23546
rect 81276 23492 81332 23494
rect 81380 23546 81436 23548
rect 81380 23494 81382 23546
rect 81382 23494 81434 23546
rect 81434 23494 81436 23546
rect 81380 23492 81436 23494
rect 81484 23546 81540 23548
rect 81484 23494 81486 23546
rect 81486 23494 81538 23546
rect 81538 23494 81540 23546
rect 81484 23492 81540 23494
rect 81116 22988 81172 23044
rect 82012 22204 82068 22260
rect 81276 21978 81332 21980
rect 81276 21926 81278 21978
rect 81278 21926 81330 21978
rect 81330 21926 81332 21978
rect 81276 21924 81332 21926
rect 81380 21978 81436 21980
rect 81380 21926 81382 21978
rect 81382 21926 81434 21978
rect 81434 21926 81436 21978
rect 81380 21924 81436 21926
rect 81484 21978 81540 21980
rect 81484 21926 81486 21978
rect 81486 21926 81538 21978
rect 81538 21926 81540 21978
rect 81484 21924 81540 21926
rect 81276 20410 81332 20412
rect 81276 20358 81278 20410
rect 81278 20358 81330 20410
rect 81330 20358 81332 20410
rect 81276 20356 81332 20358
rect 81380 20410 81436 20412
rect 81380 20358 81382 20410
rect 81382 20358 81434 20410
rect 81434 20358 81436 20410
rect 81380 20356 81436 20358
rect 81484 20410 81540 20412
rect 81484 20358 81486 20410
rect 81486 20358 81538 20410
rect 81538 20358 81540 20410
rect 81484 20356 81540 20358
rect 81004 19404 81060 19460
rect 80892 11788 80948 11844
rect 81276 18842 81332 18844
rect 81276 18790 81278 18842
rect 81278 18790 81330 18842
rect 81330 18790 81332 18842
rect 81276 18788 81332 18790
rect 81380 18842 81436 18844
rect 81380 18790 81382 18842
rect 81382 18790 81434 18842
rect 81434 18790 81436 18842
rect 81380 18788 81436 18790
rect 81484 18842 81540 18844
rect 81484 18790 81486 18842
rect 81486 18790 81538 18842
rect 81538 18790 81540 18842
rect 81484 18788 81540 18790
rect 81276 17274 81332 17276
rect 81276 17222 81278 17274
rect 81278 17222 81330 17274
rect 81330 17222 81332 17274
rect 81276 17220 81332 17222
rect 81380 17274 81436 17276
rect 81380 17222 81382 17274
rect 81382 17222 81434 17274
rect 81434 17222 81436 17274
rect 81380 17220 81436 17222
rect 81484 17274 81540 17276
rect 81484 17222 81486 17274
rect 81486 17222 81538 17274
rect 81538 17222 81540 17274
rect 81484 17220 81540 17222
rect 81276 15706 81332 15708
rect 81276 15654 81278 15706
rect 81278 15654 81330 15706
rect 81330 15654 81332 15706
rect 81276 15652 81332 15654
rect 81380 15706 81436 15708
rect 81380 15654 81382 15706
rect 81382 15654 81434 15706
rect 81434 15654 81436 15706
rect 81380 15652 81436 15654
rect 81484 15706 81540 15708
rect 81484 15654 81486 15706
rect 81486 15654 81538 15706
rect 81538 15654 81540 15706
rect 81484 15652 81540 15654
rect 81276 14138 81332 14140
rect 81276 14086 81278 14138
rect 81278 14086 81330 14138
rect 81330 14086 81332 14138
rect 81276 14084 81332 14086
rect 81380 14138 81436 14140
rect 81380 14086 81382 14138
rect 81382 14086 81434 14138
rect 81434 14086 81436 14138
rect 81380 14084 81436 14086
rect 81484 14138 81540 14140
rect 81484 14086 81486 14138
rect 81486 14086 81538 14138
rect 81538 14086 81540 14138
rect 81484 14084 81540 14086
rect 84812 20636 84868 20692
rect 82348 18620 82404 18676
rect 82012 12796 82068 12852
rect 80780 9212 80836 9268
rect 81116 12684 81172 12740
rect 80668 8540 80724 8596
rect 80780 8876 80836 8932
rect 80556 8092 80612 8148
rect 80668 8316 80724 8372
rect 81004 9826 81060 9828
rect 81004 9774 81006 9826
rect 81006 9774 81058 9826
rect 81058 9774 81060 9826
rect 81004 9772 81060 9774
rect 81004 9436 81060 9492
rect 81452 12738 81508 12740
rect 81452 12686 81454 12738
rect 81454 12686 81506 12738
rect 81506 12686 81508 12738
rect 81452 12684 81508 12686
rect 81276 12570 81332 12572
rect 81276 12518 81278 12570
rect 81278 12518 81330 12570
rect 81330 12518 81332 12570
rect 81276 12516 81332 12518
rect 81380 12570 81436 12572
rect 81380 12518 81382 12570
rect 81382 12518 81434 12570
rect 81434 12518 81436 12570
rect 81380 12516 81436 12518
rect 81484 12570 81540 12572
rect 81484 12518 81486 12570
rect 81486 12518 81538 12570
rect 81538 12518 81540 12570
rect 81484 12516 81540 12518
rect 81676 12402 81732 12404
rect 81676 12350 81678 12402
rect 81678 12350 81730 12402
rect 81730 12350 81732 12402
rect 81676 12348 81732 12350
rect 82012 12348 82068 12404
rect 82124 12908 82180 12964
rect 81340 11788 81396 11844
rect 83020 13468 83076 13524
rect 83020 13074 83076 13076
rect 83020 13022 83022 13074
rect 83022 13022 83074 13074
rect 83074 13022 83076 13074
rect 83020 13020 83076 13022
rect 82572 12402 82628 12404
rect 82572 12350 82574 12402
rect 82574 12350 82626 12402
rect 82626 12350 82628 12402
rect 82572 12348 82628 12350
rect 82236 12066 82292 12068
rect 82236 12014 82238 12066
rect 82238 12014 82290 12066
rect 82290 12014 82292 12066
rect 82236 12012 82292 12014
rect 82348 11788 82404 11844
rect 81276 11002 81332 11004
rect 81276 10950 81278 11002
rect 81278 10950 81330 11002
rect 81330 10950 81332 11002
rect 81276 10948 81332 10950
rect 81380 11002 81436 11004
rect 81380 10950 81382 11002
rect 81382 10950 81434 11002
rect 81434 10950 81436 11002
rect 81380 10948 81436 10950
rect 81484 11002 81540 11004
rect 81484 10950 81486 11002
rect 81486 10950 81538 11002
rect 81538 10950 81540 11002
rect 81484 10948 81540 10950
rect 81228 10498 81284 10500
rect 81228 10446 81230 10498
rect 81230 10446 81282 10498
rect 81282 10446 81284 10498
rect 81228 10444 81284 10446
rect 81676 9996 81732 10052
rect 81452 9826 81508 9828
rect 81452 9774 81454 9826
rect 81454 9774 81506 9826
rect 81506 9774 81508 9826
rect 81452 9772 81508 9774
rect 81788 9772 81844 9828
rect 81276 9434 81332 9436
rect 81276 9382 81278 9434
rect 81278 9382 81330 9434
rect 81330 9382 81332 9434
rect 81276 9380 81332 9382
rect 81380 9434 81436 9436
rect 81380 9382 81382 9434
rect 81382 9382 81434 9434
rect 81434 9382 81436 9434
rect 81380 9380 81436 9382
rect 81484 9434 81540 9436
rect 81484 9382 81486 9434
rect 81486 9382 81538 9434
rect 81538 9382 81540 9434
rect 81484 9380 81540 9382
rect 81564 9266 81620 9268
rect 81564 9214 81566 9266
rect 81566 9214 81618 9266
rect 81618 9214 81620 9266
rect 81564 9212 81620 9214
rect 82124 11452 82180 11508
rect 82236 10444 82292 10500
rect 82236 9826 82292 9828
rect 82236 9774 82238 9826
rect 82238 9774 82290 9826
rect 82290 9774 82292 9826
rect 82236 9772 82292 9774
rect 83244 11788 83300 11844
rect 82796 11506 82852 11508
rect 82796 11454 82798 11506
rect 82798 11454 82850 11506
rect 82850 11454 82852 11506
rect 82796 11452 82852 11454
rect 82684 10668 82740 10724
rect 82684 10444 82740 10500
rect 82348 9548 82404 9604
rect 82572 9436 82628 9492
rect 80892 8258 80948 8260
rect 80892 8206 80894 8258
rect 80894 8206 80946 8258
rect 80946 8206 80948 8258
rect 80892 8204 80948 8206
rect 80780 7644 80836 7700
rect 81004 7420 81060 7476
rect 81900 8652 81956 8708
rect 81788 8428 81844 8484
rect 81676 8316 81732 8372
rect 81340 8146 81396 8148
rect 81340 8094 81342 8146
rect 81342 8094 81394 8146
rect 81394 8094 81396 8146
rect 81340 8092 81396 8094
rect 81276 7866 81332 7868
rect 81276 7814 81278 7866
rect 81278 7814 81330 7866
rect 81330 7814 81332 7866
rect 81276 7812 81332 7814
rect 81380 7866 81436 7868
rect 81380 7814 81382 7866
rect 81382 7814 81434 7866
rect 81434 7814 81436 7866
rect 81380 7812 81436 7814
rect 81484 7866 81540 7868
rect 81484 7814 81486 7866
rect 81486 7814 81538 7866
rect 81538 7814 81540 7866
rect 81484 7812 81540 7814
rect 81564 7644 81620 7700
rect 81676 7532 81732 7588
rect 81228 7420 81284 7476
rect 80332 5906 80388 5908
rect 80332 5854 80334 5906
rect 80334 5854 80386 5906
rect 80386 5854 80388 5906
rect 80332 5852 80388 5854
rect 80444 6524 80500 6580
rect 81676 7250 81732 7252
rect 81676 7198 81678 7250
rect 81678 7198 81730 7250
rect 81730 7198 81732 7250
rect 81676 7196 81732 7198
rect 81228 6748 81284 6804
rect 81452 6578 81508 6580
rect 81452 6526 81454 6578
rect 81454 6526 81506 6578
rect 81506 6526 81508 6578
rect 81452 6524 81508 6526
rect 80780 6188 80836 6244
rect 79324 4844 79380 4900
rect 77980 4226 78036 4228
rect 77980 4174 77982 4226
rect 77982 4174 78034 4226
rect 78034 4174 78036 4226
rect 77980 4172 78036 4174
rect 79324 3724 79380 3780
rect 77644 3388 77700 3444
rect 78764 3442 78820 3444
rect 78764 3390 78766 3442
rect 78766 3390 78818 3442
rect 78818 3390 78820 3442
rect 78764 3388 78820 3390
rect 80220 5010 80276 5012
rect 80220 4958 80222 5010
rect 80222 4958 80274 5010
rect 80274 4958 80276 5010
rect 80220 4956 80276 4958
rect 80108 4898 80164 4900
rect 80108 4846 80110 4898
rect 80110 4846 80162 4898
rect 80162 4846 80164 4898
rect 80108 4844 80164 4846
rect 79996 3724 80052 3780
rect 80668 5906 80724 5908
rect 80668 5854 80670 5906
rect 80670 5854 80722 5906
rect 80722 5854 80724 5906
rect 80668 5852 80724 5854
rect 80892 5740 80948 5796
rect 81276 6298 81332 6300
rect 81276 6246 81278 6298
rect 81278 6246 81330 6298
rect 81330 6246 81332 6298
rect 81276 6244 81332 6246
rect 81380 6298 81436 6300
rect 81380 6246 81382 6298
rect 81382 6246 81434 6298
rect 81434 6246 81436 6298
rect 81380 6244 81436 6246
rect 81484 6298 81540 6300
rect 81484 6246 81486 6298
rect 81486 6246 81538 6298
rect 81538 6246 81540 6298
rect 81484 6244 81540 6246
rect 81452 6130 81508 6132
rect 81452 6078 81454 6130
rect 81454 6078 81506 6130
rect 81506 6078 81508 6130
rect 81452 6076 81508 6078
rect 81340 6018 81396 6020
rect 81340 5966 81342 6018
rect 81342 5966 81394 6018
rect 81394 5966 81396 6018
rect 81340 5964 81396 5966
rect 81228 5234 81284 5236
rect 81228 5182 81230 5234
rect 81230 5182 81282 5234
rect 81282 5182 81284 5234
rect 81228 5180 81284 5182
rect 82124 8818 82180 8820
rect 82124 8766 82126 8818
rect 82126 8766 82178 8818
rect 82178 8766 82180 8818
rect 82124 8764 82180 8766
rect 82012 8204 82068 8260
rect 82124 8316 82180 8372
rect 81116 5010 81172 5012
rect 81116 4958 81118 5010
rect 81118 4958 81170 5010
rect 81170 4958 81172 5010
rect 81116 4956 81172 4958
rect 81276 4730 81332 4732
rect 81276 4678 81278 4730
rect 81278 4678 81330 4730
rect 81330 4678 81332 4730
rect 81276 4676 81332 4678
rect 81380 4730 81436 4732
rect 81380 4678 81382 4730
rect 81382 4678 81434 4730
rect 81434 4678 81436 4730
rect 81380 4676 81436 4678
rect 81484 4730 81540 4732
rect 81484 4678 81486 4730
rect 81486 4678 81538 4730
rect 81538 4678 81540 4730
rect 81484 4676 81540 4678
rect 80444 3948 80500 4004
rect 82572 9212 82628 9268
rect 82348 7474 82404 7476
rect 82348 7422 82350 7474
rect 82350 7422 82402 7474
rect 82402 7422 82404 7474
rect 82348 7420 82404 7422
rect 82572 8652 82628 8708
rect 82124 7084 82180 7140
rect 82236 6860 82292 6916
rect 82348 6412 82404 6468
rect 82124 5906 82180 5908
rect 82124 5854 82126 5906
rect 82126 5854 82178 5906
rect 82178 5854 82180 5906
rect 82124 5852 82180 5854
rect 82236 6300 82292 6356
rect 79884 1596 79940 1652
rect 81276 3162 81332 3164
rect 81276 3110 81278 3162
rect 81278 3110 81330 3162
rect 81330 3110 81332 3162
rect 81276 3108 81332 3110
rect 81380 3162 81436 3164
rect 81380 3110 81382 3162
rect 81382 3110 81434 3162
rect 81434 3110 81436 3162
rect 81380 3108 81436 3110
rect 81484 3162 81540 3164
rect 81484 3110 81486 3162
rect 81486 3110 81538 3162
rect 81538 3110 81540 3162
rect 81484 3108 81540 3110
rect 82460 6188 82516 6244
rect 82684 6300 82740 6356
rect 82348 6130 82404 6132
rect 82348 6078 82350 6130
rect 82350 6078 82402 6130
rect 82402 6078 82404 6130
rect 82348 6076 82404 6078
rect 82572 6130 82628 6132
rect 82572 6078 82574 6130
rect 82574 6078 82626 6130
rect 82626 6078 82628 6130
rect 82572 6076 82628 6078
rect 82908 9548 82964 9604
rect 83132 9602 83188 9604
rect 83132 9550 83134 9602
rect 83134 9550 83186 9602
rect 83186 9550 83188 9602
rect 83132 9548 83188 9550
rect 83020 9042 83076 9044
rect 83020 8990 83022 9042
rect 83022 8990 83074 9042
rect 83074 8990 83076 9042
rect 83020 8988 83076 8990
rect 83468 11452 83524 11508
rect 83580 10050 83636 10052
rect 83580 9998 83582 10050
rect 83582 9998 83634 10050
rect 83634 9998 83636 10050
rect 83580 9996 83636 9998
rect 82908 6300 82964 6356
rect 83020 6972 83076 7028
rect 82684 5964 82740 6020
rect 82236 4508 82292 4564
rect 82348 4450 82404 4452
rect 82348 4398 82350 4450
rect 82350 4398 82402 4450
rect 82402 4398 82404 4450
rect 82348 4396 82404 4398
rect 82684 5292 82740 5348
rect 83132 6076 83188 6132
rect 83692 9436 83748 9492
rect 83580 8930 83636 8932
rect 83580 8878 83582 8930
rect 83582 8878 83634 8930
rect 83634 8878 83636 8930
rect 83580 8876 83636 8878
rect 83692 8370 83748 8372
rect 83692 8318 83694 8370
rect 83694 8318 83746 8370
rect 83746 8318 83748 8370
rect 83692 8316 83748 8318
rect 83468 7420 83524 7476
rect 83244 5852 83300 5908
rect 83468 6300 83524 6356
rect 83020 5740 83076 5796
rect 83468 6076 83524 6132
rect 83020 5292 83076 5348
rect 82908 4284 82964 4340
rect 83580 5404 83636 5460
rect 83468 5010 83524 5012
rect 83468 4958 83470 5010
rect 83470 4958 83522 5010
rect 83522 4958 83524 5010
rect 83468 4956 83524 4958
rect 83356 4898 83412 4900
rect 83356 4846 83358 4898
rect 83358 4846 83410 4898
rect 83410 4846 83412 4898
rect 83356 4844 83412 4846
rect 83356 4508 83412 4564
rect 86940 19180 86996 19236
rect 85932 18620 85988 18676
rect 84476 11170 84532 11172
rect 84476 11118 84478 11170
rect 84478 11118 84530 11170
rect 84530 11118 84532 11170
rect 84476 11116 84532 11118
rect 85372 13020 85428 13076
rect 84252 8764 84308 8820
rect 84028 7420 84084 7476
rect 83916 7308 83972 7364
rect 84028 7196 84084 7252
rect 83916 6524 83972 6580
rect 84140 6466 84196 6468
rect 84140 6414 84142 6466
rect 84142 6414 84194 6466
rect 84194 6414 84196 6466
rect 84140 6412 84196 6414
rect 84140 5516 84196 5572
rect 85260 9996 85316 10052
rect 86380 10892 86436 10948
rect 84588 9938 84644 9940
rect 84588 9886 84590 9938
rect 84590 9886 84642 9938
rect 84642 9886 84644 9938
rect 84588 9884 84644 9886
rect 84924 9660 84980 9716
rect 84812 8316 84868 8372
rect 84700 8092 84756 8148
rect 84252 5404 84308 5460
rect 84476 5292 84532 5348
rect 84588 6412 84644 6468
rect 84588 4956 84644 5012
rect 84028 4898 84084 4900
rect 84028 4846 84030 4898
rect 84030 4846 84082 4898
rect 84082 4846 84084 4898
rect 84028 4844 84084 4846
rect 83804 4508 83860 4564
rect 84476 4732 84532 4788
rect 84700 5404 84756 5460
rect 84252 4396 84308 4452
rect 83804 4338 83860 4340
rect 83804 4286 83806 4338
rect 83806 4286 83858 4338
rect 83858 4286 83860 4338
rect 83804 4284 83860 4286
rect 82012 1260 82068 1316
rect 85148 9548 85204 9604
rect 85036 8540 85092 8596
rect 85036 8092 85092 8148
rect 84924 4844 84980 4900
rect 85036 5852 85092 5908
rect 84812 4396 84868 4452
rect 83804 2380 83860 2436
rect 84364 3388 84420 3444
rect 85260 7980 85316 8036
rect 85260 6690 85316 6692
rect 85260 6638 85262 6690
rect 85262 6638 85314 6690
rect 85314 6638 85316 6690
rect 85260 6636 85316 6638
rect 85148 5516 85204 5572
rect 85148 4562 85204 4564
rect 85148 4510 85150 4562
rect 85150 4510 85202 4562
rect 85202 4510 85204 4562
rect 85148 4508 85204 4510
rect 85484 10332 85540 10388
rect 85484 8258 85540 8260
rect 85484 8206 85486 8258
rect 85486 8206 85538 8258
rect 85538 8206 85540 8258
rect 85484 8204 85540 8206
rect 85484 6466 85540 6468
rect 85484 6414 85486 6466
rect 85486 6414 85538 6466
rect 85538 6414 85540 6466
rect 85484 6412 85540 6414
rect 85708 9100 85764 9156
rect 85820 9996 85876 10052
rect 86156 9436 86212 9492
rect 85820 8316 85876 8372
rect 86268 8370 86324 8372
rect 86268 8318 86270 8370
rect 86270 8318 86322 8370
rect 86322 8318 86324 8370
rect 86268 8316 86324 8318
rect 86492 9042 86548 9044
rect 86492 8990 86494 9042
rect 86494 8990 86546 9042
rect 86546 8990 86548 9042
rect 86492 8988 86548 8990
rect 86492 8092 86548 8148
rect 85820 6578 85876 6580
rect 85820 6526 85822 6578
rect 85822 6526 85874 6578
rect 85874 6526 85876 6578
rect 85820 6524 85876 6526
rect 85596 6188 85652 6244
rect 87052 17724 87108 17780
rect 88844 17612 88900 17668
rect 87836 15372 87892 15428
rect 87612 10892 87668 10948
rect 86940 8316 86996 8372
rect 86828 8204 86884 8260
rect 86716 8146 86772 8148
rect 86716 8094 86718 8146
rect 86718 8094 86770 8146
rect 86770 8094 86772 8146
rect 86716 8092 86772 8094
rect 86380 6748 86436 6804
rect 85484 5964 85540 6020
rect 85484 5180 85540 5236
rect 85596 4732 85652 4788
rect 85596 4338 85652 4340
rect 85596 4286 85598 4338
rect 85598 4286 85650 4338
rect 85650 4286 85652 4338
rect 85596 4284 85652 4286
rect 85148 3442 85204 3444
rect 85148 3390 85150 3442
rect 85150 3390 85202 3442
rect 85202 3390 85204 3442
rect 85148 3388 85204 3390
rect 84812 1484 84868 1540
rect 86044 6018 86100 6020
rect 86044 5966 86046 6018
rect 86046 5966 86098 6018
rect 86098 5966 86100 6018
rect 86044 5964 86100 5966
rect 85820 4898 85876 4900
rect 85820 4846 85822 4898
rect 85822 4846 85874 4898
rect 85874 4846 85876 4898
rect 85820 4844 85876 4846
rect 86940 7980 86996 8036
rect 86716 6636 86772 6692
rect 86492 5740 86548 5796
rect 87612 10668 87668 10724
rect 87612 10108 87668 10164
rect 87500 9996 87556 10052
rect 87612 9714 87668 9716
rect 87612 9662 87614 9714
rect 87614 9662 87666 9714
rect 87666 9662 87668 9714
rect 87612 9660 87668 9662
rect 87500 9436 87556 9492
rect 87276 8258 87332 8260
rect 87276 8206 87278 8258
rect 87278 8206 87330 8258
rect 87330 8206 87332 8258
rect 87276 8204 87332 8206
rect 87052 6524 87108 6580
rect 86828 6188 86884 6244
rect 86604 5404 86660 5460
rect 87276 6748 87332 6804
rect 87500 8092 87556 8148
rect 87500 6636 87556 6692
rect 87836 8146 87892 8148
rect 87836 8094 87838 8146
rect 87838 8094 87890 8146
rect 87890 8094 87892 8146
rect 87836 8092 87892 8094
rect 87724 7532 87780 7588
rect 87724 7362 87780 7364
rect 87724 7310 87726 7362
rect 87726 7310 87778 7362
rect 87778 7310 87780 7362
rect 87724 7308 87780 7310
rect 87836 6412 87892 6468
rect 86604 4898 86660 4900
rect 86604 4846 86606 4898
rect 86606 4846 86658 4898
rect 86658 4846 86660 4898
rect 86604 4844 86660 4846
rect 85708 1036 85764 1092
rect 88396 11116 88452 11172
rect 88284 10498 88340 10500
rect 88284 10446 88286 10498
rect 88286 10446 88338 10498
rect 88338 10446 88340 10498
rect 88284 10444 88340 10446
rect 88172 9996 88228 10052
rect 88284 10108 88340 10164
rect 88172 9100 88228 9156
rect 88508 8930 88564 8932
rect 88508 8878 88510 8930
rect 88510 8878 88562 8930
rect 88562 8878 88564 8930
rect 88508 8876 88564 8878
rect 88172 6412 88228 6468
rect 87948 5180 88004 5236
rect 87612 924 87668 980
rect 88172 5234 88228 5236
rect 88172 5182 88174 5234
rect 88174 5182 88226 5234
rect 88226 5182 88228 5234
rect 88172 5180 88228 5182
rect 88508 7362 88564 7364
rect 88508 7310 88510 7362
rect 88510 7310 88562 7362
rect 88562 7310 88564 7362
rect 88508 7308 88564 7310
rect 88396 6300 88452 6356
rect 88732 7308 88788 7364
rect 88620 5068 88676 5124
rect 88732 6188 88788 6244
rect 88396 4508 88452 4564
rect 89852 16044 89908 16100
rect 89516 12124 89572 12180
rect 88956 11394 89012 11396
rect 88956 11342 88958 11394
rect 88958 11342 89010 11394
rect 89010 11342 89012 11394
rect 88956 11340 89012 11342
rect 88956 10108 89012 10164
rect 89068 9714 89124 9716
rect 89068 9662 89070 9714
rect 89070 9662 89122 9714
rect 89122 9662 89124 9714
rect 89068 9660 89124 9662
rect 89292 8092 89348 8148
rect 89628 8540 89684 8596
rect 89516 8204 89572 8260
rect 89404 8034 89460 8036
rect 89404 7982 89406 8034
rect 89406 7982 89458 8034
rect 89458 7982 89460 8034
rect 89404 7980 89460 7982
rect 90188 11900 90244 11956
rect 90412 11676 90468 11732
rect 90412 11452 90468 11508
rect 91084 11676 91140 11732
rect 91084 10556 91140 10612
rect 96636 24330 96692 24332
rect 96636 24278 96638 24330
rect 96638 24278 96690 24330
rect 96690 24278 96692 24330
rect 96636 24276 96692 24278
rect 96740 24330 96796 24332
rect 96740 24278 96742 24330
rect 96742 24278 96794 24330
rect 96794 24278 96796 24330
rect 96740 24276 96796 24278
rect 96844 24330 96900 24332
rect 96844 24278 96846 24330
rect 96846 24278 96898 24330
rect 96898 24278 96900 24330
rect 96844 24276 96900 24278
rect 96636 22762 96692 22764
rect 96636 22710 96638 22762
rect 96638 22710 96690 22762
rect 96690 22710 96692 22762
rect 96636 22708 96692 22710
rect 96740 22762 96796 22764
rect 96740 22710 96742 22762
rect 96742 22710 96794 22762
rect 96794 22710 96796 22762
rect 96740 22708 96796 22710
rect 96844 22762 96900 22764
rect 96844 22710 96846 22762
rect 96846 22710 96898 22762
rect 96898 22710 96900 22762
rect 96844 22708 96900 22710
rect 96636 21194 96692 21196
rect 96636 21142 96638 21194
rect 96638 21142 96690 21194
rect 96690 21142 96692 21194
rect 96636 21140 96692 21142
rect 96740 21194 96796 21196
rect 96740 21142 96742 21194
rect 96742 21142 96794 21194
rect 96794 21142 96796 21194
rect 96740 21140 96796 21142
rect 96844 21194 96900 21196
rect 96844 21142 96846 21194
rect 96846 21142 96898 21194
rect 96898 21142 96900 21194
rect 96844 21140 96900 21142
rect 100716 24444 100772 24500
rect 99036 20860 99092 20916
rect 96636 19626 96692 19628
rect 96636 19574 96638 19626
rect 96638 19574 96690 19626
rect 96690 19574 96692 19626
rect 96636 19572 96692 19574
rect 96740 19626 96796 19628
rect 96740 19574 96742 19626
rect 96742 19574 96794 19626
rect 96794 19574 96796 19626
rect 96740 19572 96796 19574
rect 96844 19626 96900 19628
rect 96844 19574 96846 19626
rect 96846 19574 96898 19626
rect 96898 19574 96900 19626
rect 96844 19572 96900 19574
rect 94444 19068 94500 19124
rect 92204 17836 92260 17892
rect 91532 11788 91588 11844
rect 91756 13804 91812 13860
rect 91644 10498 91700 10500
rect 91644 10446 91646 10498
rect 91646 10446 91698 10498
rect 91698 10446 91700 10498
rect 91644 10444 91700 10446
rect 90188 9266 90244 9268
rect 90188 9214 90190 9266
rect 90190 9214 90242 9266
rect 90242 9214 90244 9266
rect 90188 9212 90244 9214
rect 90300 8540 90356 8596
rect 90188 8258 90244 8260
rect 90188 8206 90190 8258
rect 90190 8206 90242 8258
rect 90242 8206 90244 8258
rect 90188 8204 90244 8206
rect 89852 7980 89908 8036
rect 88956 6300 89012 6356
rect 89180 6188 89236 6244
rect 89068 5964 89124 6020
rect 89740 7196 89796 7252
rect 90860 7980 90916 8036
rect 90748 7532 90804 7588
rect 90188 7196 90244 7252
rect 89852 6748 89908 6804
rect 90076 6188 90132 6244
rect 88844 4508 88900 4564
rect 89180 4060 89236 4116
rect 89292 5292 89348 5348
rect 89740 5010 89796 5012
rect 89740 4958 89742 5010
rect 89742 4958 89794 5010
rect 89794 4958 89796 5010
rect 89740 4956 89796 4958
rect 90524 6466 90580 6468
rect 90524 6414 90526 6466
rect 90526 6414 90578 6466
rect 90578 6414 90580 6466
rect 90524 6412 90580 6414
rect 90636 6188 90692 6244
rect 90972 5964 91028 6020
rect 90748 5906 90804 5908
rect 90748 5854 90750 5906
rect 90750 5854 90802 5906
rect 90802 5854 90804 5906
rect 90748 5852 90804 5854
rect 90972 5794 91028 5796
rect 90972 5742 90974 5794
rect 90974 5742 91026 5794
rect 91026 5742 91028 5794
rect 90972 5740 91028 5742
rect 91308 7980 91364 8036
rect 89964 4844 90020 4900
rect 90188 4844 90244 4900
rect 90076 4562 90132 4564
rect 90076 4510 90078 4562
rect 90078 4510 90130 4562
rect 90130 4510 90132 4562
rect 90076 4508 90132 4510
rect 88060 3500 88116 3556
rect 89404 4338 89460 4340
rect 89404 4286 89406 4338
rect 89406 4286 89458 4338
rect 89458 4286 89460 4338
rect 89404 4284 89460 4286
rect 90412 5180 90468 5236
rect 91084 5068 91140 5124
rect 90972 5010 91028 5012
rect 90972 4958 90974 5010
rect 90974 4958 91026 5010
rect 91026 4958 91028 5010
rect 90972 4956 91028 4958
rect 90524 4898 90580 4900
rect 90524 4846 90526 4898
rect 90526 4846 90578 4898
rect 90578 4846 90580 4898
rect 90524 4844 90580 4846
rect 91308 5234 91364 5236
rect 91308 5182 91310 5234
rect 91310 5182 91362 5234
rect 91362 5182 91364 5234
rect 91308 5180 91364 5182
rect 91644 8316 91700 8372
rect 92092 12236 92148 12292
rect 91868 8540 91924 8596
rect 91980 8146 92036 8148
rect 91980 8094 91982 8146
rect 91982 8094 92034 8146
rect 92034 8094 92036 8146
rect 91980 8092 92036 8094
rect 91532 6690 91588 6692
rect 91532 6638 91534 6690
rect 91534 6638 91586 6690
rect 91586 6638 91588 6690
rect 91532 6636 91588 6638
rect 91868 6300 91924 6356
rect 91644 6018 91700 6020
rect 91644 5966 91646 6018
rect 91646 5966 91698 6018
rect 91698 5966 91700 6018
rect 91644 5964 91700 5966
rect 91980 5852 92036 5908
rect 91532 5740 91588 5796
rect 91756 5794 91812 5796
rect 91756 5742 91758 5794
rect 91758 5742 91810 5794
rect 91810 5742 91812 5794
rect 91756 5740 91812 5742
rect 91868 5516 91924 5572
rect 91644 5404 91700 5460
rect 91308 4732 91364 4788
rect 91644 4732 91700 4788
rect 90972 4226 91028 4228
rect 90972 4174 90974 4226
rect 90974 4174 91026 4226
rect 91026 4174 91028 4226
rect 90972 4172 91028 4174
rect 91756 4060 91812 4116
rect 89628 3554 89684 3556
rect 89628 3502 89630 3554
rect 89630 3502 89682 3554
rect 89682 3502 89684 3554
rect 89628 3500 89684 3502
rect 89292 1372 89348 1428
rect 89404 3388 89460 3444
rect 90524 3442 90580 3444
rect 90524 3390 90526 3442
rect 90526 3390 90578 3442
rect 90578 3390 90580 3442
rect 90524 3388 90580 3390
rect 91084 3388 91140 3444
rect 92092 5292 92148 5348
rect 91980 3948 92036 4004
rect 93436 15484 93492 15540
rect 92316 15372 92372 15428
rect 92428 11394 92484 11396
rect 92428 11342 92430 11394
rect 92430 11342 92482 11394
rect 92482 11342 92484 11394
rect 92428 11340 92484 11342
rect 93212 8876 93268 8932
rect 92428 8540 92484 8596
rect 92988 8428 93044 8484
rect 92428 8370 92484 8372
rect 92428 8318 92430 8370
rect 92430 8318 92482 8370
rect 92482 8318 92484 8370
rect 92428 8316 92484 8318
rect 93100 8092 93156 8148
rect 93212 7196 93268 7252
rect 93996 14700 94052 14756
rect 93660 12124 93716 12180
rect 92540 6188 92596 6244
rect 93548 11788 93604 11844
rect 93548 7698 93604 7700
rect 93548 7646 93550 7698
rect 93550 7646 93602 7698
rect 93602 7646 93604 7698
rect 93548 7644 93604 7646
rect 93100 6300 93156 6356
rect 92316 5180 92372 5236
rect 92428 4508 92484 4564
rect 93212 5010 93268 5012
rect 93212 4958 93214 5010
rect 93214 4958 93266 5010
rect 93266 4958 93268 5010
rect 93212 4956 93268 4958
rect 92540 4284 92596 4340
rect 93772 11394 93828 11396
rect 93772 11342 93774 11394
rect 93774 11342 93826 11394
rect 93826 11342 93828 11394
rect 93772 11340 93828 11342
rect 94108 13916 94164 13972
rect 95564 19068 95620 19124
rect 95228 16268 95284 16324
rect 94780 16156 94836 16212
rect 94220 11340 94276 11396
rect 93996 9660 94052 9716
rect 93772 8428 93828 8484
rect 94220 9100 94276 9156
rect 94108 8428 94164 8484
rect 94220 8370 94276 8372
rect 94220 8318 94222 8370
rect 94222 8318 94274 8370
rect 94274 8318 94276 8370
rect 94220 8316 94276 8318
rect 95116 10444 95172 10500
rect 95004 9602 95060 9604
rect 95004 9550 95006 9602
rect 95006 9550 95058 9602
rect 95058 9550 95060 9602
rect 95004 9548 95060 9550
rect 95340 10220 95396 10276
rect 96636 18058 96692 18060
rect 96636 18006 96638 18058
rect 96638 18006 96690 18058
rect 96690 18006 96692 18058
rect 96636 18004 96692 18006
rect 96740 18058 96796 18060
rect 96740 18006 96742 18058
rect 96742 18006 96794 18058
rect 96794 18006 96796 18058
rect 96740 18004 96796 18006
rect 96844 18058 96900 18060
rect 96844 18006 96846 18058
rect 96846 18006 96898 18058
rect 96898 18006 96900 18058
rect 96844 18004 96900 18006
rect 95564 9996 95620 10052
rect 95676 17388 95732 17444
rect 94780 8482 94836 8484
rect 94780 8430 94782 8482
rect 94782 8430 94834 8482
rect 94834 8430 94836 8482
rect 94780 8428 94836 8430
rect 95228 8428 95284 8484
rect 94556 8092 94612 8148
rect 94780 7980 94836 8036
rect 94444 7698 94500 7700
rect 94444 7646 94446 7698
rect 94446 7646 94498 7698
rect 94498 7646 94500 7698
rect 94444 7644 94500 7646
rect 93996 7532 94052 7588
rect 93660 5404 93716 5460
rect 93772 7420 93828 7476
rect 93772 6076 93828 6132
rect 94892 7868 94948 7924
rect 95004 8092 95060 8148
rect 95340 8370 95396 8372
rect 95340 8318 95342 8370
rect 95342 8318 95394 8370
rect 95394 8318 95396 8370
rect 95340 8316 95396 8318
rect 97580 16828 97636 16884
rect 96636 16490 96692 16492
rect 96636 16438 96638 16490
rect 96638 16438 96690 16490
rect 96690 16438 96692 16490
rect 96636 16436 96692 16438
rect 96740 16490 96796 16492
rect 96740 16438 96742 16490
rect 96742 16438 96794 16490
rect 96794 16438 96796 16490
rect 96740 16436 96796 16438
rect 96844 16490 96900 16492
rect 96844 16438 96846 16490
rect 96846 16438 96898 16490
rect 96898 16438 96900 16490
rect 96844 16436 96900 16438
rect 96348 15932 96404 15988
rect 97132 15820 97188 15876
rect 96012 11116 96068 11172
rect 96012 10220 96068 10276
rect 95788 8316 95844 8372
rect 95452 8204 95508 8260
rect 95564 7980 95620 8036
rect 95228 7756 95284 7812
rect 95340 7644 95396 7700
rect 95228 7586 95284 7588
rect 95228 7534 95230 7586
rect 95230 7534 95282 7586
rect 95282 7534 95284 7586
rect 95228 7532 95284 7534
rect 95676 7586 95732 7588
rect 95676 7534 95678 7586
rect 95678 7534 95730 7586
rect 95730 7534 95732 7586
rect 95676 7532 95732 7534
rect 95228 6860 95284 6916
rect 95116 6636 95172 6692
rect 96636 14922 96692 14924
rect 96636 14870 96638 14922
rect 96638 14870 96690 14922
rect 96690 14870 96692 14922
rect 96636 14868 96692 14870
rect 96740 14922 96796 14924
rect 96740 14870 96742 14922
rect 96742 14870 96794 14922
rect 96794 14870 96796 14922
rect 96740 14868 96796 14870
rect 96844 14922 96900 14924
rect 96844 14870 96846 14922
rect 96846 14870 96898 14922
rect 96898 14870 96900 14922
rect 96844 14868 96900 14870
rect 96636 13354 96692 13356
rect 96636 13302 96638 13354
rect 96638 13302 96690 13354
rect 96690 13302 96692 13354
rect 96636 13300 96692 13302
rect 96740 13354 96796 13356
rect 96740 13302 96742 13354
rect 96742 13302 96794 13354
rect 96794 13302 96796 13354
rect 96740 13300 96796 13302
rect 96844 13354 96900 13356
rect 96844 13302 96846 13354
rect 96846 13302 96898 13354
rect 96898 13302 96900 13354
rect 96844 13300 96900 13302
rect 96636 11786 96692 11788
rect 96636 11734 96638 11786
rect 96638 11734 96690 11786
rect 96690 11734 96692 11786
rect 96636 11732 96692 11734
rect 96740 11786 96796 11788
rect 96740 11734 96742 11786
rect 96742 11734 96794 11786
rect 96794 11734 96796 11786
rect 96740 11732 96796 11734
rect 96844 11786 96900 11788
rect 96844 11734 96846 11786
rect 96846 11734 96898 11786
rect 96898 11734 96900 11786
rect 96844 11732 96900 11734
rect 97132 11676 97188 11732
rect 97692 11676 97748 11732
rect 96460 11340 96516 11396
rect 96636 10218 96692 10220
rect 96636 10166 96638 10218
rect 96638 10166 96690 10218
rect 96690 10166 96692 10218
rect 96636 10164 96692 10166
rect 96740 10218 96796 10220
rect 96740 10166 96742 10218
rect 96742 10166 96794 10218
rect 96794 10166 96796 10218
rect 96740 10164 96796 10166
rect 96844 10218 96900 10220
rect 96844 10166 96846 10218
rect 96846 10166 96898 10218
rect 96898 10166 96900 10218
rect 96844 10164 96900 10166
rect 96572 9714 96628 9716
rect 96572 9662 96574 9714
rect 96574 9662 96626 9714
rect 96626 9662 96628 9714
rect 96572 9660 96628 9662
rect 98140 11676 98196 11732
rect 98140 11340 98196 11396
rect 97244 10498 97300 10500
rect 97244 10446 97246 10498
rect 97246 10446 97298 10498
rect 97298 10446 97300 10498
rect 97244 10444 97300 10446
rect 97804 10444 97860 10500
rect 98252 10892 98308 10948
rect 96236 9266 96292 9268
rect 96236 9214 96238 9266
rect 96238 9214 96290 9266
rect 96290 9214 96292 9266
rect 96236 9212 96292 9214
rect 96348 8258 96404 8260
rect 96348 8206 96350 8258
rect 96350 8206 96402 8258
rect 96402 8206 96404 8258
rect 96348 8204 96404 8206
rect 96572 8818 96628 8820
rect 96572 8766 96574 8818
rect 96574 8766 96626 8818
rect 96626 8766 96628 8818
rect 96572 8764 96628 8766
rect 96636 8650 96692 8652
rect 96636 8598 96638 8650
rect 96638 8598 96690 8650
rect 96690 8598 96692 8650
rect 96636 8596 96692 8598
rect 96740 8650 96796 8652
rect 96740 8598 96742 8650
rect 96742 8598 96794 8650
rect 96794 8598 96796 8650
rect 96740 8596 96796 8598
rect 96844 8650 96900 8652
rect 96844 8598 96846 8650
rect 96846 8598 96898 8650
rect 96898 8598 96900 8650
rect 96844 8596 96900 8598
rect 96684 8316 96740 8372
rect 96236 8034 96292 8036
rect 96236 7982 96238 8034
rect 96238 7982 96290 8034
rect 96290 7982 96292 8034
rect 96236 7980 96292 7982
rect 96460 7868 96516 7924
rect 97468 9548 97524 9604
rect 97020 7644 97076 7700
rect 96124 7362 96180 7364
rect 96124 7310 96126 7362
rect 96126 7310 96178 7362
rect 96178 7310 96180 7362
rect 96124 7308 96180 7310
rect 95900 6690 95956 6692
rect 95900 6638 95902 6690
rect 95902 6638 95954 6690
rect 95954 6638 95956 6690
rect 95900 6636 95956 6638
rect 94556 6300 94612 6356
rect 95564 6300 95620 6356
rect 95004 6188 95060 6244
rect 93772 5068 93828 5124
rect 93660 4956 93716 5012
rect 94108 5010 94164 5012
rect 94108 4958 94110 5010
rect 94110 4958 94162 5010
rect 94162 4958 94164 5010
rect 94108 4956 94164 4958
rect 93324 4562 93380 4564
rect 93324 4510 93326 4562
rect 93326 4510 93378 4562
rect 93378 4510 93380 4562
rect 93324 4508 93380 4510
rect 92204 4172 92260 4228
rect 92988 4396 93044 4452
rect 92764 4338 92820 4340
rect 92764 4286 92766 4338
rect 92766 4286 92818 4338
rect 92818 4286 92820 4338
rect 92764 4284 92820 4286
rect 92652 3724 92708 3780
rect 92764 3500 92820 3556
rect 91868 2380 91924 2436
rect 92876 3442 92932 3444
rect 92876 3390 92878 3442
rect 92878 3390 92930 3442
rect 92930 3390 92932 3442
rect 92876 3388 92932 3390
rect 93772 4226 93828 4228
rect 93772 4174 93774 4226
rect 93774 4174 93826 4226
rect 93826 4174 93828 4226
rect 93772 4172 93828 4174
rect 95004 5180 95060 5236
rect 94668 4844 94724 4900
rect 94108 3164 94164 3220
rect 94444 3724 94500 3780
rect 93324 2716 93380 2772
rect 95340 4898 95396 4900
rect 95340 4846 95342 4898
rect 95342 4846 95394 4898
rect 95394 4846 95396 4898
rect 95340 4844 95396 4846
rect 95116 4508 95172 4564
rect 96236 6860 96292 6916
rect 96236 6690 96292 6692
rect 96236 6638 96238 6690
rect 96238 6638 96290 6690
rect 96290 6638 96292 6690
rect 96236 6636 96292 6638
rect 97132 9100 97188 9156
rect 96636 7082 96692 7084
rect 96636 7030 96638 7082
rect 96638 7030 96690 7082
rect 96690 7030 96692 7082
rect 96636 7028 96692 7030
rect 96740 7082 96796 7084
rect 96740 7030 96742 7082
rect 96742 7030 96794 7082
rect 96794 7030 96796 7082
rect 96740 7028 96796 7030
rect 96844 7082 96900 7084
rect 96844 7030 96846 7082
rect 96846 7030 96898 7082
rect 96898 7030 96900 7082
rect 96844 7028 96900 7030
rect 96684 6860 96740 6916
rect 96236 6018 96292 6020
rect 96236 5966 96238 6018
rect 96238 5966 96290 6018
rect 96290 5966 96292 6018
rect 96236 5964 96292 5966
rect 96012 5682 96068 5684
rect 96012 5630 96014 5682
rect 96014 5630 96066 5682
rect 96066 5630 96068 5682
rect 96012 5628 96068 5630
rect 96636 5514 96692 5516
rect 96636 5462 96638 5514
rect 96638 5462 96690 5514
rect 96690 5462 96692 5514
rect 96636 5460 96692 5462
rect 96740 5514 96796 5516
rect 96740 5462 96742 5514
rect 96742 5462 96794 5514
rect 96794 5462 96796 5514
rect 96740 5460 96796 5462
rect 96844 5514 96900 5516
rect 96844 5462 96846 5514
rect 96846 5462 96898 5514
rect 96898 5462 96900 5514
rect 96844 5460 96900 5462
rect 96348 5068 96404 5124
rect 96124 5010 96180 5012
rect 96124 4958 96126 5010
rect 96126 4958 96178 5010
rect 96178 4958 96180 5010
rect 96124 4956 96180 4958
rect 95340 3724 95396 3780
rect 94780 3612 94836 3668
rect 94668 3554 94724 3556
rect 94668 3502 94670 3554
rect 94670 3502 94722 3554
rect 94722 3502 94724 3554
rect 94668 3500 94724 3502
rect 96124 3388 96180 3444
rect 96796 4956 96852 5012
rect 96348 4396 96404 4452
rect 96460 4844 96516 4900
rect 96796 4396 96852 4452
rect 97356 9154 97412 9156
rect 97356 9102 97358 9154
rect 97358 9102 97410 9154
rect 97410 9102 97412 9154
rect 97356 9100 97412 9102
rect 97244 8316 97300 8372
rect 97244 7644 97300 7700
rect 97356 7868 97412 7924
rect 97580 9212 97636 9268
rect 97692 9548 97748 9604
rect 98364 9714 98420 9716
rect 98364 9662 98366 9714
rect 98366 9662 98418 9714
rect 98418 9662 98420 9714
rect 98364 9660 98420 9662
rect 97804 9324 97860 9380
rect 98364 9436 98420 9492
rect 97580 7868 97636 7924
rect 97804 7868 97860 7924
rect 97692 7756 97748 7812
rect 97244 7362 97300 7364
rect 97244 7310 97246 7362
rect 97246 7310 97298 7362
rect 97298 7310 97300 7362
rect 97244 7308 97300 7310
rect 97580 7196 97636 7252
rect 97244 6972 97300 7028
rect 97468 6690 97524 6692
rect 97468 6638 97470 6690
rect 97470 6638 97522 6690
rect 97522 6638 97524 6690
rect 97468 6636 97524 6638
rect 97356 5964 97412 6020
rect 97132 5180 97188 5236
rect 97020 4898 97076 4900
rect 97020 4846 97022 4898
rect 97022 4846 97074 4898
rect 97074 4846 97076 4898
rect 97020 4844 97076 4846
rect 97692 6748 97748 6804
rect 98252 9100 98308 9156
rect 98028 7644 98084 7700
rect 98140 7532 98196 7588
rect 98140 7196 98196 7252
rect 98252 7868 98308 7924
rect 98252 7084 98308 7140
rect 97020 4508 97076 4564
rect 97356 4450 97412 4452
rect 97356 4398 97358 4450
rect 97358 4398 97410 4450
rect 97410 4398 97412 4450
rect 97356 4396 97412 4398
rect 96908 4060 96964 4116
rect 96636 3946 96692 3948
rect 96636 3894 96638 3946
rect 96638 3894 96690 3946
rect 96690 3894 96692 3946
rect 96636 3892 96692 3894
rect 96740 3946 96796 3948
rect 96740 3894 96742 3946
rect 96742 3894 96794 3946
rect 96794 3894 96796 3946
rect 96740 3892 96796 3894
rect 96844 3946 96900 3948
rect 96844 3894 96846 3946
rect 96846 3894 96898 3946
rect 96898 3894 96900 3946
rect 96844 3892 96900 3894
rect 97244 3442 97300 3444
rect 97244 3390 97246 3442
rect 97246 3390 97298 3442
rect 97298 3390 97300 3442
rect 97244 3388 97300 3390
rect 96236 3276 96292 3332
rect 98812 11676 98868 11732
rect 100604 14476 100660 14532
rect 100492 13916 100548 13972
rect 100380 12738 100436 12740
rect 100380 12686 100382 12738
rect 100382 12686 100434 12738
rect 100434 12686 100436 12738
rect 100380 12684 100436 12686
rect 100156 11676 100212 11732
rect 99148 11170 99204 11172
rect 99148 11118 99150 11170
rect 99150 11118 99202 11170
rect 99202 11118 99204 11170
rect 99148 11116 99204 11118
rect 99036 10892 99092 10948
rect 98700 10108 98756 10164
rect 98812 9660 98868 9716
rect 99148 9826 99204 9828
rect 99148 9774 99150 9826
rect 99150 9774 99202 9826
rect 99202 9774 99204 9826
rect 99148 9772 99204 9774
rect 99148 9324 99204 9380
rect 98588 7420 98644 7476
rect 98700 7362 98756 7364
rect 98700 7310 98702 7362
rect 98702 7310 98754 7362
rect 98754 7310 98756 7362
rect 98700 7308 98756 7310
rect 98588 6748 98644 6804
rect 99372 9602 99428 9604
rect 99372 9550 99374 9602
rect 99374 9550 99426 9602
rect 99426 9550 99428 9602
rect 99372 9548 99428 9550
rect 99484 9154 99540 9156
rect 99484 9102 99486 9154
rect 99486 9102 99538 9154
rect 99538 9102 99540 9154
rect 99484 9100 99540 9102
rect 99148 8258 99204 8260
rect 99148 8206 99150 8258
rect 99150 8206 99202 8258
rect 99202 8206 99204 8258
rect 99148 8204 99204 8206
rect 99260 8092 99316 8148
rect 99148 7362 99204 7364
rect 99148 7310 99150 7362
rect 99150 7310 99202 7362
rect 99202 7310 99204 7362
rect 99148 7308 99204 7310
rect 99260 6860 99316 6916
rect 99036 6578 99092 6580
rect 99036 6526 99038 6578
rect 99038 6526 99090 6578
rect 99090 6526 99092 6578
rect 99036 6524 99092 6526
rect 98924 5906 98980 5908
rect 98924 5854 98926 5906
rect 98926 5854 98978 5906
rect 98978 5854 98980 5906
rect 98924 5852 98980 5854
rect 98924 5180 98980 5236
rect 98812 5068 98868 5124
rect 98812 4844 98868 4900
rect 99932 11282 99988 11284
rect 99932 11230 99934 11282
rect 99934 11230 99986 11282
rect 99986 11230 99988 11282
rect 99932 11228 99988 11230
rect 100044 11004 100100 11060
rect 99820 9602 99876 9604
rect 99820 9550 99822 9602
rect 99822 9550 99874 9602
rect 99874 9550 99876 9602
rect 99820 9548 99876 9550
rect 99932 9100 99988 9156
rect 99708 8764 99764 8820
rect 100156 10610 100212 10612
rect 100156 10558 100158 10610
rect 100158 10558 100210 10610
rect 100210 10558 100212 10610
rect 100156 10556 100212 10558
rect 100268 11900 100324 11956
rect 100380 10892 100436 10948
rect 100716 11116 100772 11172
rect 102396 30268 102452 30324
rect 102060 21420 102116 21476
rect 101276 18956 101332 19012
rect 101164 12684 101220 12740
rect 101052 11340 101108 11396
rect 101164 11170 101220 11172
rect 101164 11118 101166 11170
rect 101166 11118 101218 11170
rect 101218 11118 101220 11170
rect 101164 11116 101220 11118
rect 100268 9772 100324 9828
rect 100380 9548 100436 9604
rect 99708 8204 99764 8260
rect 99820 8146 99876 8148
rect 99820 8094 99822 8146
rect 99822 8094 99874 8146
rect 99874 8094 99876 8146
rect 99820 8092 99876 8094
rect 99596 7756 99652 7812
rect 99484 6690 99540 6692
rect 99484 6638 99486 6690
rect 99486 6638 99538 6690
rect 99538 6638 99540 6690
rect 99484 6636 99540 6638
rect 99708 7698 99764 7700
rect 99708 7646 99710 7698
rect 99710 7646 99762 7698
rect 99762 7646 99764 7698
rect 99708 7644 99764 7646
rect 100156 8370 100212 8372
rect 100156 8318 100158 8370
rect 100158 8318 100210 8370
rect 100210 8318 100212 8370
rect 100156 8316 100212 8318
rect 100156 7980 100212 8036
rect 100156 6860 100212 6916
rect 99932 6690 99988 6692
rect 99932 6638 99934 6690
rect 99934 6638 99986 6690
rect 99986 6638 99988 6690
rect 99932 6636 99988 6638
rect 98476 4620 98532 4676
rect 99820 5234 99876 5236
rect 99820 5182 99822 5234
rect 99822 5182 99874 5234
rect 99874 5182 99876 5234
rect 99820 5180 99876 5182
rect 97692 1596 97748 1652
rect 97804 4172 97860 4228
rect 98700 4226 98756 4228
rect 98700 4174 98702 4226
rect 98702 4174 98754 4226
rect 98754 4174 98756 4226
rect 98700 4172 98756 4174
rect 98924 4060 98980 4116
rect 98476 3554 98532 3556
rect 98476 3502 98478 3554
rect 98478 3502 98530 3554
rect 98530 3502 98532 3554
rect 98476 3500 98532 3502
rect 100604 9100 100660 9156
rect 100492 8652 100548 8708
rect 100604 8204 100660 8260
rect 100492 7756 100548 7812
rect 100492 7474 100548 7476
rect 100492 7422 100494 7474
rect 100494 7422 100546 7474
rect 100546 7422 100548 7474
rect 100492 7420 100548 7422
rect 100380 7308 100436 7364
rect 100268 5404 100324 5460
rect 100380 4956 100436 5012
rect 100268 4620 100324 4676
rect 99484 3388 99540 3444
rect 98140 3330 98196 3332
rect 98140 3278 98142 3330
rect 98142 3278 98194 3330
rect 98194 3278 98196 3330
rect 98140 3276 98196 3278
rect 98588 1596 98644 1652
rect 100044 3276 100100 3332
rect 100940 9548 100996 9604
rect 100940 9266 100996 9268
rect 100940 9214 100942 9266
rect 100942 9214 100994 9266
rect 100994 9214 100996 9266
rect 100940 9212 100996 9214
rect 100828 7980 100884 8036
rect 100940 7698 100996 7700
rect 100940 7646 100942 7698
rect 100942 7646 100994 7698
rect 100994 7646 100996 7698
rect 100940 7644 100996 7646
rect 101052 7420 101108 7476
rect 100716 5628 100772 5684
rect 101724 11340 101780 11396
rect 101500 11004 101556 11060
rect 101276 9548 101332 9604
rect 101388 8988 101444 9044
rect 101164 5964 101220 6020
rect 101052 5234 101108 5236
rect 101052 5182 101054 5234
rect 101054 5182 101106 5234
rect 101106 5182 101108 5234
rect 101052 5180 101108 5182
rect 101276 8428 101332 8484
rect 101388 8258 101444 8260
rect 101388 8206 101390 8258
rect 101390 8206 101442 8258
rect 101442 8206 101444 8258
rect 101388 8204 101444 8206
rect 101612 8652 101668 8708
rect 101612 8146 101668 8148
rect 101612 8094 101614 8146
rect 101614 8094 101666 8146
rect 101666 8094 101668 8146
rect 101612 8092 101668 8094
rect 101500 7868 101556 7924
rect 101500 7698 101556 7700
rect 101500 7646 101502 7698
rect 101502 7646 101554 7698
rect 101554 7646 101556 7698
rect 101500 7644 101556 7646
rect 104412 25452 104468 25508
rect 104300 21308 104356 21364
rect 104076 11900 104132 11956
rect 104300 11452 104356 11508
rect 101836 6524 101892 6580
rect 101276 4844 101332 4900
rect 101612 6300 101668 6356
rect 102508 11228 102564 11284
rect 102732 10220 102788 10276
rect 103628 10780 103684 10836
rect 103516 10722 103572 10724
rect 103516 10670 103518 10722
rect 103518 10670 103570 10722
rect 103570 10670 103572 10722
rect 103516 10668 103572 10670
rect 102844 8988 102900 9044
rect 102956 10498 103012 10500
rect 102956 10446 102958 10498
rect 102958 10446 103010 10498
rect 103010 10446 103012 10498
rect 102956 10444 103012 10446
rect 103292 10220 103348 10276
rect 102396 8428 102452 8484
rect 103068 10108 103124 10164
rect 102396 8034 102452 8036
rect 102396 7982 102398 8034
rect 102398 7982 102450 8034
rect 102450 7982 102452 8034
rect 102396 7980 102452 7982
rect 104188 10722 104244 10724
rect 104188 10670 104190 10722
rect 104190 10670 104242 10722
rect 104242 10670 104244 10722
rect 104188 10668 104244 10670
rect 107660 116450 107716 116452
rect 107660 116398 107662 116450
rect 107662 116398 107714 116450
rect 107714 116398 107716 116450
rect 107660 116396 107716 116398
rect 108332 116562 108388 116564
rect 108332 116510 108334 116562
rect 108334 116510 108386 116562
rect 108386 116510 108388 116562
rect 108332 116508 108388 116510
rect 115836 116620 115892 116676
rect 116732 116620 116788 116676
rect 111996 116058 112052 116060
rect 111996 116006 111998 116058
rect 111998 116006 112050 116058
rect 112050 116006 112052 116058
rect 111996 116004 112052 116006
rect 112100 116058 112156 116060
rect 112100 116006 112102 116058
rect 112102 116006 112154 116058
rect 112154 116006 112156 116058
rect 112100 116004 112156 116006
rect 112204 116058 112260 116060
rect 112204 116006 112206 116058
rect 112206 116006 112258 116058
rect 112258 116006 112260 116058
rect 112204 116004 112260 116006
rect 107996 115724 108052 115780
rect 108556 115778 108612 115780
rect 108556 115726 108558 115778
rect 108558 115726 108610 115778
rect 108610 115726 108612 115778
rect 108556 115724 108612 115726
rect 110460 115612 110516 115668
rect 106092 23772 106148 23828
rect 105756 14588 105812 14644
rect 105420 12012 105476 12068
rect 104076 10332 104132 10388
rect 103964 10220 104020 10276
rect 102956 7868 103012 7924
rect 102732 7474 102788 7476
rect 102732 7422 102734 7474
rect 102734 7422 102786 7474
rect 102786 7422 102788 7474
rect 102732 7420 102788 7422
rect 102284 6300 102340 6356
rect 101836 6018 101892 6020
rect 101836 5966 101838 6018
rect 101838 5966 101890 6018
rect 101890 5966 101892 6018
rect 101836 5964 101892 5966
rect 101724 5292 101780 5348
rect 101500 4396 101556 4452
rect 102396 6972 102452 7028
rect 102060 5346 102116 5348
rect 102060 5294 102062 5346
rect 102062 5294 102114 5346
rect 102114 5294 102116 5346
rect 102060 5292 102116 5294
rect 102508 6748 102564 6804
rect 102396 5292 102452 5348
rect 102620 6524 102676 6580
rect 102844 4956 102900 5012
rect 103516 7980 103572 8036
rect 103628 7420 103684 7476
rect 103068 6300 103124 6356
rect 103292 5292 103348 5348
rect 102956 4844 103012 4900
rect 103292 4844 103348 4900
rect 104300 9042 104356 9044
rect 104300 8990 104302 9042
rect 104302 8990 104354 9042
rect 104354 8990 104356 9042
rect 104300 8988 104356 8990
rect 104748 11452 104804 11508
rect 104524 8876 104580 8932
rect 104412 8258 104468 8260
rect 104412 8206 104414 8258
rect 104414 8206 104466 8258
rect 104466 8206 104468 8258
rect 104412 8204 104468 8206
rect 104188 7586 104244 7588
rect 104188 7534 104190 7586
rect 104190 7534 104242 7586
rect 104242 7534 104244 7586
rect 104188 7532 104244 7534
rect 104188 7196 104244 7252
rect 103964 6860 104020 6916
rect 104188 6690 104244 6692
rect 104188 6638 104190 6690
rect 104190 6638 104242 6690
rect 104242 6638 104244 6690
rect 104188 6636 104244 6638
rect 103852 6300 103908 6356
rect 104076 5516 104132 5572
rect 103740 5122 103796 5124
rect 103740 5070 103742 5122
rect 103742 5070 103794 5122
rect 103794 5070 103796 5122
rect 103740 5068 103796 5070
rect 102172 4508 102228 4564
rect 100716 3442 100772 3444
rect 100716 3390 100718 3442
rect 100718 3390 100770 3442
rect 100770 3390 100772 3442
rect 100716 3388 100772 3390
rect 101164 3388 101220 3444
rect 100492 1372 100548 1428
rect 102172 4338 102228 4340
rect 102172 4286 102174 4338
rect 102174 4286 102226 4338
rect 102226 4286 102228 4338
rect 102172 4284 102228 4286
rect 102396 3724 102452 3780
rect 103292 4450 103348 4452
rect 103292 4398 103294 4450
rect 103294 4398 103346 4450
rect 103346 4398 103348 4450
rect 103292 4396 103348 4398
rect 104188 4338 104244 4340
rect 104188 4286 104190 4338
rect 104190 4286 104242 4338
rect 104242 4286 104244 4338
rect 104188 4284 104244 4286
rect 104412 6636 104468 6692
rect 104524 6578 104580 6580
rect 104524 6526 104526 6578
rect 104526 6526 104578 6578
rect 104578 6526 104580 6578
rect 104524 6524 104580 6526
rect 104412 6300 104468 6356
rect 104412 4956 104468 5012
rect 104524 4732 104580 4788
rect 105980 12066 106036 12068
rect 105980 12014 105982 12066
rect 105982 12014 106034 12066
rect 106034 12014 106036 12066
rect 105980 12012 106036 12014
rect 105756 10780 105812 10836
rect 105308 10722 105364 10724
rect 105308 10670 105310 10722
rect 105310 10670 105362 10722
rect 105362 10670 105364 10722
rect 105308 10668 105364 10670
rect 105532 10108 105588 10164
rect 108668 27132 108724 27188
rect 107100 18508 107156 18564
rect 106876 14028 106932 14084
rect 106764 12012 106820 12068
rect 106428 10834 106484 10836
rect 106428 10782 106430 10834
rect 106430 10782 106482 10834
rect 106482 10782 106484 10834
rect 106428 10780 106484 10782
rect 105196 8876 105252 8932
rect 105196 8540 105252 8596
rect 104860 8204 104916 8260
rect 105084 8034 105140 8036
rect 105084 7982 105086 8034
rect 105086 7982 105138 8034
rect 105138 7982 105140 8034
rect 105084 7980 105140 7982
rect 105084 6690 105140 6692
rect 105084 6638 105086 6690
rect 105086 6638 105138 6690
rect 105138 6638 105140 6690
rect 105084 6636 105140 6638
rect 105308 6636 105364 6692
rect 106092 10108 106148 10164
rect 106428 10332 106484 10388
rect 106652 10332 106708 10388
rect 105980 9602 106036 9604
rect 105980 9550 105982 9602
rect 105982 9550 106034 9602
rect 106034 9550 106036 9602
rect 105980 9548 106036 9550
rect 105532 8876 105588 8932
rect 105532 8204 105588 8260
rect 105644 8764 105700 8820
rect 105980 8540 106036 8596
rect 106092 8428 106148 8484
rect 105756 8034 105812 8036
rect 105756 7982 105758 8034
rect 105758 7982 105810 8034
rect 105810 7982 105812 8034
rect 105756 7980 105812 7982
rect 105532 7698 105588 7700
rect 105532 7646 105534 7698
rect 105534 7646 105586 7698
rect 105586 7646 105588 7698
rect 105532 7644 105588 7646
rect 105756 7532 105812 7588
rect 105644 6578 105700 6580
rect 105644 6526 105646 6578
rect 105646 6526 105698 6578
rect 105698 6526 105700 6578
rect 105644 6524 105700 6526
rect 104972 5852 105028 5908
rect 104748 4396 104804 4452
rect 101948 3442 102004 3444
rect 101948 3390 101950 3442
rect 101950 3390 102002 3442
rect 102002 3390 102004 3442
rect 101948 3388 102004 3390
rect 104076 3442 104132 3444
rect 104076 3390 104078 3442
rect 104078 3390 104130 3442
rect 104130 3390 104132 3442
rect 104076 3388 104132 3390
rect 104524 3388 104580 3444
rect 101836 3276 101892 3332
rect 102844 3276 102900 3332
rect 104748 3612 104804 3668
rect 104636 3276 104692 3332
rect 105196 5516 105252 5572
rect 105644 6076 105700 6132
rect 105420 5794 105476 5796
rect 105420 5742 105422 5794
rect 105422 5742 105474 5794
rect 105474 5742 105476 5794
rect 105420 5740 105476 5742
rect 105644 5628 105700 5684
rect 105644 5292 105700 5348
rect 105420 5180 105476 5236
rect 105308 4732 105364 4788
rect 106204 7532 106260 7588
rect 106428 7474 106484 7476
rect 106428 7422 106430 7474
rect 106430 7422 106482 7474
rect 106482 7422 106484 7474
rect 106428 7420 106484 7422
rect 105868 6524 105924 6580
rect 105980 6412 106036 6468
rect 106092 6636 106148 6692
rect 105868 5068 105924 5124
rect 105980 4844 106036 4900
rect 106652 8034 106708 8036
rect 106652 7982 106654 8034
rect 106654 7982 106706 8034
rect 106706 7982 106708 8034
rect 106652 7980 106708 7982
rect 106316 5234 106372 5236
rect 106316 5182 106318 5234
rect 106318 5182 106370 5234
rect 106370 5182 106372 5234
rect 106316 5180 106372 5182
rect 105308 4562 105364 4564
rect 105308 4510 105310 4562
rect 105310 4510 105362 4562
rect 105362 4510 105364 4562
rect 105308 4508 105364 4510
rect 106540 5740 106596 5796
rect 106652 7084 106708 7140
rect 106988 10332 107044 10388
rect 106876 8092 106932 8148
rect 107212 12684 107268 12740
rect 106876 7868 106932 7924
rect 106764 6690 106820 6692
rect 106764 6638 106766 6690
rect 106766 6638 106818 6690
rect 106818 6638 106820 6690
rect 106764 6636 106820 6638
rect 106652 5404 106708 5460
rect 106876 6076 106932 6132
rect 106428 4508 106484 4564
rect 106540 4956 106596 5012
rect 105420 4284 105476 4340
rect 105980 4338 106036 4340
rect 105980 4286 105982 4338
rect 105982 4286 106034 4338
rect 106034 4286 106036 4338
rect 105980 4284 106036 4286
rect 106204 4172 106260 4228
rect 105084 2156 105140 2212
rect 106428 3442 106484 3444
rect 106428 3390 106430 3442
rect 106430 3390 106482 3442
rect 106482 3390 106484 3442
rect 106428 3388 106484 3390
rect 108108 12066 108164 12068
rect 108108 12014 108110 12066
rect 108110 12014 108162 12066
rect 108162 12014 108164 12066
rect 108108 12012 108164 12014
rect 107884 10556 107940 10612
rect 107100 7644 107156 7700
rect 107100 6972 107156 7028
rect 107212 8146 107268 8148
rect 107212 8094 107214 8146
rect 107214 8094 107266 8146
rect 107266 8094 107268 8146
rect 107212 8092 107268 8094
rect 107212 6748 107268 6804
rect 107100 6636 107156 6692
rect 108332 10556 108388 10612
rect 107884 8988 107940 9044
rect 108108 8764 108164 8820
rect 107436 7698 107492 7700
rect 107436 7646 107438 7698
rect 107438 7646 107490 7698
rect 107490 7646 107492 7698
rect 107436 7644 107492 7646
rect 107324 6636 107380 6692
rect 107100 6018 107156 6020
rect 107100 5966 107102 6018
rect 107102 5966 107154 6018
rect 107154 5966 107156 6018
rect 107100 5964 107156 5966
rect 107436 5964 107492 6020
rect 107436 5740 107492 5796
rect 107324 4732 107380 4788
rect 107996 8034 108052 8036
rect 107996 7982 107998 8034
rect 107998 7982 108050 8034
rect 108050 7982 108052 8034
rect 107996 7980 108052 7982
rect 107884 7868 107940 7924
rect 107660 7756 107716 7812
rect 107660 5516 107716 5572
rect 107996 7586 108052 7588
rect 107996 7534 107998 7586
rect 107998 7534 108050 7586
rect 108050 7534 108052 7586
rect 107996 7532 108052 7534
rect 107996 6972 108052 7028
rect 108668 10332 108724 10388
rect 108556 10220 108612 10276
rect 108668 9100 108724 9156
rect 108444 8316 108500 8372
rect 107996 5852 108052 5908
rect 107548 4844 107604 4900
rect 107100 4226 107156 4228
rect 107100 4174 107102 4226
rect 107102 4174 107154 4226
rect 107154 4174 107156 4226
rect 107100 4172 107156 4174
rect 108220 7084 108276 7140
rect 108220 6300 108276 6356
rect 108108 4284 108164 4340
rect 107548 4172 107604 4228
rect 107548 3554 107604 3556
rect 107548 3502 107550 3554
rect 107550 3502 107602 3554
rect 107602 3502 107604 3554
rect 107548 3500 107604 3502
rect 108332 5010 108388 5012
rect 108332 4958 108334 5010
rect 108334 4958 108386 5010
rect 108386 4958 108388 5010
rect 108332 4956 108388 4958
rect 108556 7644 108612 7700
rect 108556 6860 108612 6916
rect 110796 115666 110852 115668
rect 110796 115614 110798 115666
rect 110798 115614 110850 115666
rect 110850 115614 110852 115666
rect 110796 115612 110852 115614
rect 113036 115554 113092 115556
rect 113036 115502 113038 115554
rect 113038 115502 113090 115554
rect 113090 115502 113092 115554
rect 113036 115500 113092 115502
rect 113932 115500 113988 115556
rect 111996 114490 112052 114492
rect 111996 114438 111998 114490
rect 111998 114438 112050 114490
rect 112050 114438 112052 114490
rect 111996 114436 112052 114438
rect 112100 114490 112156 114492
rect 112100 114438 112102 114490
rect 112102 114438 112154 114490
rect 112154 114438 112156 114490
rect 112100 114436 112156 114438
rect 112204 114490 112260 114492
rect 112204 114438 112206 114490
rect 112206 114438 112258 114490
rect 112258 114438 112260 114490
rect 112204 114436 112260 114438
rect 111996 112922 112052 112924
rect 111996 112870 111998 112922
rect 111998 112870 112050 112922
rect 112050 112870 112052 112922
rect 111996 112868 112052 112870
rect 112100 112922 112156 112924
rect 112100 112870 112102 112922
rect 112102 112870 112154 112922
rect 112154 112870 112156 112922
rect 112100 112868 112156 112870
rect 112204 112922 112260 112924
rect 112204 112870 112206 112922
rect 112206 112870 112258 112922
rect 112258 112870 112260 112922
rect 112204 112868 112260 112870
rect 111996 111354 112052 111356
rect 111996 111302 111998 111354
rect 111998 111302 112050 111354
rect 112050 111302 112052 111354
rect 111996 111300 112052 111302
rect 112100 111354 112156 111356
rect 112100 111302 112102 111354
rect 112102 111302 112154 111354
rect 112154 111302 112156 111354
rect 112100 111300 112156 111302
rect 112204 111354 112260 111356
rect 112204 111302 112206 111354
rect 112206 111302 112258 111354
rect 112258 111302 112260 111354
rect 112204 111300 112260 111302
rect 111996 109786 112052 109788
rect 111996 109734 111998 109786
rect 111998 109734 112050 109786
rect 112050 109734 112052 109786
rect 111996 109732 112052 109734
rect 112100 109786 112156 109788
rect 112100 109734 112102 109786
rect 112102 109734 112154 109786
rect 112154 109734 112156 109786
rect 112100 109732 112156 109734
rect 112204 109786 112260 109788
rect 112204 109734 112206 109786
rect 112206 109734 112258 109786
rect 112258 109734 112260 109786
rect 112204 109732 112260 109734
rect 111996 108218 112052 108220
rect 111996 108166 111998 108218
rect 111998 108166 112050 108218
rect 112050 108166 112052 108218
rect 111996 108164 112052 108166
rect 112100 108218 112156 108220
rect 112100 108166 112102 108218
rect 112102 108166 112154 108218
rect 112154 108166 112156 108218
rect 112100 108164 112156 108166
rect 112204 108218 112260 108220
rect 112204 108166 112206 108218
rect 112206 108166 112258 108218
rect 112258 108166 112260 108218
rect 112204 108164 112260 108166
rect 111996 106650 112052 106652
rect 111996 106598 111998 106650
rect 111998 106598 112050 106650
rect 112050 106598 112052 106650
rect 111996 106596 112052 106598
rect 112100 106650 112156 106652
rect 112100 106598 112102 106650
rect 112102 106598 112154 106650
rect 112154 106598 112156 106650
rect 112100 106596 112156 106598
rect 112204 106650 112260 106652
rect 112204 106598 112206 106650
rect 112206 106598 112258 106650
rect 112258 106598 112260 106650
rect 112204 106596 112260 106598
rect 111996 105082 112052 105084
rect 111996 105030 111998 105082
rect 111998 105030 112050 105082
rect 112050 105030 112052 105082
rect 111996 105028 112052 105030
rect 112100 105082 112156 105084
rect 112100 105030 112102 105082
rect 112102 105030 112154 105082
rect 112154 105030 112156 105082
rect 112100 105028 112156 105030
rect 112204 105082 112260 105084
rect 112204 105030 112206 105082
rect 112206 105030 112258 105082
rect 112258 105030 112260 105082
rect 112204 105028 112260 105030
rect 111996 103514 112052 103516
rect 111996 103462 111998 103514
rect 111998 103462 112050 103514
rect 112050 103462 112052 103514
rect 111996 103460 112052 103462
rect 112100 103514 112156 103516
rect 112100 103462 112102 103514
rect 112102 103462 112154 103514
rect 112154 103462 112156 103514
rect 112100 103460 112156 103462
rect 112204 103514 112260 103516
rect 112204 103462 112206 103514
rect 112206 103462 112258 103514
rect 112258 103462 112260 103514
rect 112204 103460 112260 103462
rect 111996 101946 112052 101948
rect 111996 101894 111998 101946
rect 111998 101894 112050 101946
rect 112050 101894 112052 101946
rect 111996 101892 112052 101894
rect 112100 101946 112156 101948
rect 112100 101894 112102 101946
rect 112102 101894 112154 101946
rect 112154 101894 112156 101946
rect 112100 101892 112156 101894
rect 112204 101946 112260 101948
rect 112204 101894 112206 101946
rect 112206 101894 112258 101946
rect 112258 101894 112260 101946
rect 112204 101892 112260 101894
rect 111996 100378 112052 100380
rect 111996 100326 111998 100378
rect 111998 100326 112050 100378
rect 112050 100326 112052 100378
rect 111996 100324 112052 100326
rect 112100 100378 112156 100380
rect 112100 100326 112102 100378
rect 112102 100326 112154 100378
rect 112154 100326 112156 100378
rect 112100 100324 112156 100326
rect 112204 100378 112260 100380
rect 112204 100326 112206 100378
rect 112206 100326 112258 100378
rect 112258 100326 112260 100378
rect 112204 100324 112260 100326
rect 111996 98810 112052 98812
rect 111996 98758 111998 98810
rect 111998 98758 112050 98810
rect 112050 98758 112052 98810
rect 111996 98756 112052 98758
rect 112100 98810 112156 98812
rect 112100 98758 112102 98810
rect 112102 98758 112154 98810
rect 112154 98758 112156 98810
rect 112100 98756 112156 98758
rect 112204 98810 112260 98812
rect 112204 98758 112206 98810
rect 112206 98758 112258 98810
rect 112258 98758 112260 98810
rect 112204 98756 112260 98758
rect 111996 97242 112052 97244
rect 111996 97190 111998 97242
rect 111998 97190 112050 97242
rect 112050 97190 112052 97242
rect 111996 97188 112052 97190
rect 112100 97242 112156 97244
rect 112100 97190 112102 97242
rect 112102 97190 112154 97242
rect 112154 97190 112156 97242
rect 112100 97188 112156 97190
rect 112204 97242 112260 97244
rect 112204 97190 112206 97242
rect 112206 97190 112258 97242
rect 112258 97190 112260 97242
rect 112204 97188 112260 97190
rect 111996 95674 112052 95676
rect 111996 95622 111998 95674
rect 111998 95622 112050 95674
rect 112050 95622 112052 95674
rect 111996 95620 112052 95622
rect 112100 95674 112156 95676
rect 112100 95622 112102 95674
rect 112102 95622 112154 95674
rect 112154 95622 112156 95674
rect 112100 95620 112156 95622
rect 112204 95674 112260 95676
rect 112204 95622 112206 95674
rect 112206 95622 112258 95674
rect 112258 95622 112260 95674
rect 112204 95620 112260 95622
rect 111996 94106 112052 94108
rect 111996 94054 111998 94106
rect 111998 94054 112050 94106
rect 112050 94054 112052 94106
rect 111996 94052 112052 94054
rect 112100 94106 112156 94108
rect 112100 94054 112102 94106
rect 112102 94054 112154 94106
rect 112154 94054 112156 94106
rect 112100 94052 112156 94054
rect 112204 94106 112260 94108
rect 112204 94054 112206 94106
rect 112206 94054 112258 94106
rect 112258 94054 112260 94106
rect 112204 94052 112260 94054
rect 111996 92538 112052 92540
rect 111996 92486 111998 92538
rect 111998 92486 112050 92538
rect 112050 92486 112052 92538
rect 111996 92484 112052 92486
rect 112100 92538 112156 92540
rect 112100 92486 112102 92538
rect 112102 92486 112154 92538
rect 112154 92486 112156 92538
rect 112100 92484 112156 92486
rect 112204 92538 112260 92540
rect 112204 92486 112206 92538
rect 112206 92486 112258 92538
rect 112258 92486 112260 92538
rect 112204 92484 112260 92486
rect 111996 90970 112052 90972
rect 111996 90918 111998 90970
rect 111998 90918 112050 90970
rect 112050 90918 112052 90970
rect 111996 90916 112052 90918
rect 112100 90970 112156 90972
rect 112100 90918 112102 90970
rect 112102 90918 112154 90970
rect 112154 90918 112156 90970
rect 112100 90916 112156 90918
rect 112204 90970 112260 90972
rect 112204 90918 112206 90970
rect 112206 90918 112258 90970
rect 112258 90918 112260 90970
rect 112204 90916 112260 90918
rect 111996 89402 112052 89404
rect 111996 89350 111998 89402
rect 111998 89350 112050 89402
rect 112050 89350 112052 89402
rect 111996 89348 112052 89350
rect 112100 89402 112156 89404
rect 112100 89350 112102 89402
rect 112102 89350 112154 89402
rect 112154 89350 112156 89402
rect 112100 89348 112156 89350
rect 112204 89402 112260 89404
rect 112204 89350 112206 89402
rect 112206 89350 112258 89402
rect 112258 89350 112260 89402
rect 112204 89348 112260 89350
rect 111996 87834 112052 87836
rect 111996 87782 111998 87834
rect 111998 87782 112050 87834
rect 112050 87782 112052 87834
rect 111996 87780 112052 87782
rect 112100 87834 112156 87836
rect 112100 87782 112102 87834
rect 112102 87782 112154 87834
rect 112154 87782 112156 87834
rect 112100 87780 112156 87782
rect 112204 87834 112260 87836
rect 112204 87782 112206 87834
rect 112206 87782 112258 87834
rect 112258 87782 112260 87834
rect 112204 87780 112260 87782
rect 111996 86266 112052 86268
rect 111996 86214 111998 86266
rect 111998 86214 112050 86266
rect 112050 86214 112052 86266
rect 111996 86212 112052 86214
rect 112100 86266 112156 86268
rect 112100 86214 112102 86266
rect 112102 86214 112154 86266
rect 112154 86214 112156 86266
rect 112100 86212 112156 86214
rect 112204 86266 112260 86268
rect 112204 86214 112206 86266
rect 112206 86214 112258 86266
rect 112258 86214 112260 86266
rect 112204 86212 112260 86214
rect 111996 84698 112052 84700
rect 111996 84646 111998 84698
rect 111998 84646 112050 84698
rect 112050 84646 112052 84698
rect 111996 84644 112052 84646
rect 112100 84698 112156 84700
rect 112100 84646 112102 84698
rect 112102 84646 112154 84698
rect 112154 84646 112156 84698
rect 112100 84644 112156 84646
rect 112204 84698 112260 84700
rect 112204 84646 112206 84698
rect 112206 84646 112258 84698
rect 112258 84646 112260 84698
rect 112204 84644 112260 84646
rect 111996 83130 112052 83132
rect 111996 83078 111998 83130
rect 111998 83078 112050 83130
rect 112050 83078 112052 83130
rect 111996 83076 112052 83078
rect 112100 83130 112156 83132
rect 112100 83078 112102 83130
rect 112102 83078 112154 83130
rect 112154 83078 112156 83130
rect 112100 83076 112156 83078
rect 112204 83130 112260 83132
rect 112204 83078 112206 83130
rect 112206 83078 112258 83130
rect 112258 83078 112260 83130
rect 112204 83076 112260 83078
rect 111996 81562 112052 81564
rect 111996 81510 111998 81562
rect 111998 81510 112050 81562
rect 112050 81510 112052 81562
rect 111996 81508 112052 81510
rect 112100 81562 112156 81564
rect 112100 81510 112102 81562
rect 112102 81510 112154 81562
rect 112154 81510 112156 81562
rect 112100 81508 112156 81510
rect 112204 81562 112260 81564
rect 112204 81510 112206 81562
rect 112206 81510 112258 81562
rect 112258 81510 112260 81562
rect 112204 81508 112260 81510
rect 111996 79994 112052 79996
rect 111996 79942 111998 79994
rect 111998 79942 112050 79994
rect 112050 79942 112052 79994
rect 111996 79940 112052 79942
rect 112100 79994 112156 79996
rect 112100 79942 112102 79994
rect 112102 79942 112154 79994
rect 112154 79942 112156 79994
rect 112100 79940 112156 79942
rect 112204 79994 112260 79996
rect 112204 79942 112206 79994
rect 112206 79942 112258 79994
rect 112258 79942 112260 79994
rect 112204 79940 112260 79942
rect 111996 78426 112052 78428
rect 111996 78374 111998 78426
rect 111998 78374 112050 78426
rect 112050 78374 112052 78426
rect 111996 78372 112052 78374
rect 112100 78426 112156 78428
rect 112100 78374 112102 78426
rect 112102 78374 112154 78426
rect 112154 78374 112156 78426
rect 112100 78372 112156 78374
rect 112204 78426 112260 78428
rect 112204 78374 112206 78426
rect 112206 78374 112258 78426
rect 112258 78374 112260 78426
rect 112204 78372 112260 78374
rect 111996 76858 112052 76860
rect 111996 76806 111998 76858
rect 111998 76806 112050 76858
rect 112050 76806 112052 76858
rect 111996 76804 112052 76806
rect 112100 76858 112156 76860
rect 112100 76806 112102 76858
rect 112102 76806 112154 76858
rect 112154 76806 112156 76858
rect 112100 76804 112156 76806
rect 112204 76858 112260 76860
rect 112204 76806 112206 76858
rect 112206 76806 112258 76858
rect 112258 76806 112260 76858
rect 112204 76804 112260 76806
rect 111996 75290 112052 75292
rect 111996 75238 111998 75290
rect 111998 75238 112050 75290
rect 112050 75238 112052 75290
rect 111996 75236 112052 75238
rect 112100 75290 112156 75292
rect 112100 75238 112102 75290
rect 112102 75238 112154 75290
rect 112154 75238 112156 75290
rect 112100 75236 112156 75238
rect 112204 75290 112260 75292
rect 112204 75238 112206 75290
rect 112206 75238 112258 75290
rect 112258 75238 112260 75290
rect 112204 75236 112260 75238
rect 111996 73722 112052 73724
rect 111996 73670 111998 73722
rect 111998 73670 112050 73722
rect 112050 73670 112052 73722
rect 111996 73668 112052 73670
rect 112100 73722 112156 73724
rect 112100 73670 112102 73722
rect 112102 73670 112154 73722
rect 112154 73670 112156 73722
rect 112100 73668 112156 73670
rect 112204 73722 112260 73724
rect 112204 73670 112206 73722
rect 112206 73670 112258 73722
rect 112258 73670 112260 73722
rect 112204 73668 112260 73670
rect 111996 72154 112052 72156
rect 111996 72102 111998 72154
rect 111998 72102 112050 72154
rect 112050 72102 112052 72154
rect 111996 72100 112052 72102
rect 112100 72154 112156 72156
rect 112100 72102 112102 72154
rect 112102 72102 112154 72154
rect 112154 72102 112156 72154
rect 112100 72100 112156 72102
rect 112204 72154 112260 72156
rect 112204 72102 112206 72154
rect 112206 72102 112258 72154
rect 112258 72102 112260 72154
rect 112204 72100 112260 72102
rect 111996 70586 112052 70588
rect 111996 70534 111998 70586
rect 111998 70534 112050 70586
rect 112050 70534 112052 70586
rect 111996 70532 112052 70534
rect 112100 70586 112156 70588
rect 112100 70534 112102 70586
rect 112102 70534 112154 70586
rect 112154 70534 112156 70586
rect 112100 70532 112156 70534
rect 112204 70586 112260 70588
rect 112204 70534 112206 70586
rect 112206 70534 112258 70586
rect 112258 70534 112260 70586
rect 112204 70532 112260 70534
rect 111996 69018 112052 69020
rect 111996 68966 111998 69018
rect 111998 68966 112050 69018
rect 112050 68966 112052 69018
rect 111996 68964 112052 68966
rect 112100 69018 112156 69020
rect 112100 68966 112102 69018
rect 112102 68966 112154 69018
rect 112154 68966 112156 69018
rect 112100 68964 112156 68966
rect 112204 69018 112260 69020
rect 112204 68966 112206 69018
rect 112206 68966 112258 69018
rect 112258 68966 112260 69018
rect 112204 68964 112260 68966
rect 111996 67450 112052 67452
rect 111996 67398 111998 67450
rect 111998 67398 112050 67450
rect 112050 67398 112052 67450
rect 111996 67396 112052 67398
rect 112100 67450 112156 67452
rect 112100 67398 112102 67450
rect 112102 67398 112154 67450
rect 112154 67398 112156 67450
rect 112100 67396 112156 67398
rect 112204 67450 112260 67452
rect 112204 67398 112206 67450
rect 112206 67398 112258 67450
rect 112258 67398 112260 67450
rect 112204 67396 112260 67398
rect 111996 65882 112052 65884
rect 111996 65830 111998 65882
rect 111998 65830 112050 65882
rect 112050 65830 112052 65882
rect 111996 65828 112052 65830
rect 112100 65882 112156 65884
rect 112100 65830 112102 65882
rect 112102 65830 112154 65882
rect 112154 65830 112156 65882
rect 112100 65828 112156 65830
rect 112204 65882 112260 65884
rect 112204 65830 112206 65882
rect 112206 65830 112258 65882
rect 112258 65830 112260 65882
rect 112204 65828 112260 65830
rect 111996 64314 112052 64316
rect 111996 64262 111998 64314
rect 111998 64262 112050 64314
rect 112050 64262 112052 64314
rect 111996 64260 112052 64262
rect 112100 64314 112156 64316
rect 112100 64262 112102 64314
rect 112102 64262 112154 64314
rect 112154 64262 112156 64314
rect 112100 64260 112156 64262
rect 112204 64314 112260 64316
rect 112204 64262 112206 64314
rect 112206 64262 112258 64314
rect 112258 64262 112260 64314
rect 112204 64260 112260 64262
rect 111996 62746 112052 62748
rect 111996 62694 111998 62746
rect 111998 62694 112050 62746
rect 112050 62694 112052 62746
rect 111996 62692 112052 62694
rect 112100 62746 112156 62748
rect 112100 62694 112102 62746
rect 112102 62694 112154 62746
rect 112154 62694 112156 62746
rect 112100 62692 112156 62694
rect 112204 62746 112260 62748
rect 112204 62694 112206 62746
rect 112206 62694 112258 62746
rect 112258 62694 112260 62746
rect 112204 62692 112260 62694
rect 111996 61178 112052 61180
rect 111996 61126 111998 61178
rect 111998 61126 112050 61178
rect 112050 61126 112052 61178
rect 111996 61124 112052 61126
rect 112100 61178 112156 61180
rect 112100 61126 112102 61178
rect 112102 61126 112154 61178
rect 112154 61126 112156 61178
rect 112100 61124 112156 61126
rect 112204 61178 112260 61180
rect 112204 61126 112206 61178
rect 112206 61126 112258 61178
rect 112258 61126 112260 61178
rect 112204 61124 112260 61126
rect 111996 59610 112052 59612
rect 111996 59558 111998 59610
rect 111998 59558 112050 59610
rect 112050 59558 112052 59610
rect 111996 59556 112052 59558
rect 112100 59610 112156 59612
rect 112100 59558 112102 59610
rect 112102 59558 112154 59610
rect 112154 59558 112156 59610
rect 112100 59556 112156 59558
rect 112204 59610 112260 59612
rect 112204 59558 112206 59610
rect 112206 59558 112258 59610
rect 112258 59558 112260 59610
rect 112204 59556 112260 59558
rect 111996 58042 112052 58044
rect 111996 57990 111998 58042
rect 111998 57990 112050 58042
rect 112050 57990 112052 58042
rect 111996 57988 112052 57990
rect 112100 58042 112156 58044
rect 112100 57990 112102 58042
rect 112102 57990 112154 58042
rect 112154 57990 112156 58042
rect 112100 57988 112156 57990
rect 112204 58042 112260 58044
rect 112204 57990 112206 58042
rect 112206 57990 112258 58042
rect 112258 57990 112260 58042
rect 112204 57988 112260 57990
rect 111996 56474 112052 56476
rect 111996 56422 111998 56474
rect 111998 56422 112050 56474
rect 112050 56422 112052 56474
rect 111996 56420 112052 56422
rect 112100 56474 112156 56476
rect 112100 56422 112102 56474
rect 112102 56422 112154 56474
rect 112154 56422 112156 56474
rect 112100 56420 112156 56422
rect 112204 56474 112260 56476
rect 112204 56422 112206 56474
rect 112206 56422 112258 56474
rect 112258 56422 112260 56474
rect 112204 56420 112260 56422
rect 111996 54906 112052 54908
rect 111996 54854 111998 54906
rect 111998 54854 112050 54906
rect 112050 54854 112052 54906
rect 111996 54852 112052 54854
rect 112100 54906 112156 54908
rect 112100 54854 112102 54906
rect 112102 54854 112154 54906
rect 112154 54854 112156 54906
rect 112100 54852 112156 54854
rect 112204 54906 112260 54908
rect 112204 54854 112206 54906
rect 112206 54854 112258 54906
rect 112258 54854 112260 54906
rect 112204 54852 112260 54854
rect 111996 53338 112052 53340
rect 111996 53286 111998 53338
rect 111998 53286 112050 53338
rect 112050 53286 112052 53338
rect 111996 53284 112052 53286
rect 112100 53338 112156 53340
rect 112100 53286 112102 53338
rect 112102 53286 112154 53338
rect 112154 53286 112156 53338
rect 112100 53284 112156 53286
rect 112204 53338 112260 53340
rect 112204 53286 112206 53338
rect 112206 53286 112258 53338
rect 112258 53286 112260 53338
rect 112204 53284 112260 53286
rect 111996 51770 112052 51772
rect 111996 51718 111998 51770
rect 111998 51718 112050 51770
rect 112050 51718 112052 51770
rect 111996 51716 112052 51718
rect 112100 51770 112156 51772
rect 112100 51718 112102 51770
rect 112102 51718 112154 51770
rect 112154 51718 112156 51770
rect 112100 51716 112156 51718
rect 112204 51770 112260 51772
rect 112204 51718 112206 51770
rect 112206 51718 112258 51770
rect 112258 51718 112260 51770
rect 112204 51716 112260 51718
rect 111996 50202 112052 50204
rect 111996 50150 111998 50202
rect 111998 50150 112050 50202
rect 112050 50150 112052 50202
rect 111996 50148 112052 50150
rect 112100 50202 112156 50204
rect 112100 50150 112102 50202
rect 112102 50150 112154 50202
rect 112154 50150 112156 50202
rect 112100 50148 112156 50150
rect 112204 50202 112260 50204
rect 112204 50150 112206 50202
rect 112206 50150 112258 50202
rect 112258 50150 112260 50202
rect 112204 50148 112260 50150
rect 111996 48634 112052 48636
rect 111996 48582 111998 48634
rect 111998 48582 112050 48634
rect 112050 48582 112052 48634
rect 111996 48580 112052 48582
rect 112100 48634 112156 48636
rect 112100 48582 112102 48634
rect 112102 48582 112154 48634
rect 112154 48582 112156 48634
rect 112100 48580 112156 48582
rect 112204 48634 112260 48636
rect 112204 48582 112206 48634
rect 112206 48582 112258 48634
rect 112258 48582 112260 48634
rect 112204 48580 112260 48582
rect 111996 47066 112052 47068
rect 111996 47014 111998 47066
rect 111998 47014 112050 47066
rect 112050 47014 112052 47066
rect 111996 47012 112052 47014
rect 112100 47066 112156 47068
rect 112100 47014 112102 47066
rect 112102 47014 112154 47066
rect 112154 47014 112156 47066
rect 112100 47012 112156 47014
rect 112204 47066 112260 47068
rect 112204 47014 112206 47066
rect 112206 47014 112258 47066
rect 112258 47014 112260 47066
rect 112204 47012 112260 47014
rect 111996 45498 112052 45500
rect 111996 45446 111998 45498
rect 111998 45446 112050 45498
rect 112050 45446 112052 45498
rect 111996 45444 112052 45446
rect 112100 45498 112156 45500
rect 112100 45446 112102 45498
rect 112102 45446 112154 45498
rect 112154 45446 112156 45498
rect 112100 45444 112156 45446
rect 112204 45498 112260 45500
rect 112204 45446 112206 45498
rect 112206 45446 112258 45498
rect 112258 45446 112260 45498
rect 112204 45444 112260 45446
rect 111996 43930 112052 43932
rect 111996 43878 111998 43930
rect 111998 43878 112050 43930
rect 112050 43878 112052 43930
rect 111996 43876 112052 43878
rect 112100 43930 112156 43932
rect 112100 43878 112102 43930
rect 112102 43878 112154 43930
rect 112154 43878 112156 43930
rect 112100 43876 112156 43878
rect 112204 43930 112260 43932
rect 112204 43878 112206 43930
rect 112206 43878 112258 43930
rect 112258 43878 112260 43930
rect 112204 43876 112260 43878
rect 111996 42362 112052 42364
rect 111996 42310 111998 42362
rect 111998 42310 112050 42362
rect 112050 42310 112052 42362
rect 111996 42308 112052 42310
rect 112100 42362 112156 42364
rect 112100 42310 112102 42362
rect 112102 42310 112154 42362
rect 112154 42310 112156 42362
rect 112100 42308 112156 42310
rect 112204 42362 112260 42364
rect 112204 42310 112206 42362
rect 112206 42310 112258 42362
rect 112258 42310 112260 42362
rect 112204 42308 112260 42310
rect 111996 40794 112052 40796
rect 111996 40742 111998 40794
rect 111998 40742 112050 40794
rect 112050 40742 112052 40794
rect 111996 40740 112052 40742
rect 112100 40794 112156 40796
rect 112100 40742 112102 40794
rect 112102 40742 112154 40794
rect 112154 40742 112156 40794
rect 112100 40740 112156 40742
rect 112204 40794 112260 40796
rect 112204 40742 112206 40794
rect 112206 40742 112258 40794
rect 112258 40742 112260 40794
rect 112204 40740 112260 40742
rect 111996 39226 112052 39228
rect 111996 39174 111998 39226
rect 111998 39174 112050 39226
rect 112050 39174 112052 39226
rect 111996 39172 112052 39174
rect 112100 39226 112156 39228
rect 112100 39174 112102 39226
rect 112102 39174 112154 39226
rect 112154 39174 112156 39226
rect 112100 39172 112156 39174
rect 112204 39226 112260 39228
rect 112204 39174 112206 39226
rect 112206 39174 112258 39226
rect 112258 39174 112260 39226
rect 112204 39172 112260 39174
rect 111996 37658 112052 37660
rect 111996 37606 111998 37658
rect 111998 37606 112050 37658
rect 112050 37606 112052 37658
rect 111996 37604 112052 37606
rect 112100 37658 112156 37660
rect 112100 37606 112102 37658
rect 112102 37606 112154 37658
rect 112154 37606 112156 37658
rect 112100 37604 112156 37606
rect 112204 37658 112260 37660
rect 112204 37606 112206 37658
rect 112206 37606 112258 37658
rect 112258 37606 112260 37658
rect 112204 37604 112260 37606
rect 111996 36090 112052 36092
rect 111996 36038 111998 36090
rect 111998 36038 112050 36090
rect 112050 36038 112052 36090
rect 111996 36036 112052 36038
rect 112100 36090 112156 36092
rect 112100 36038 112102 36090
rect 112102 36038 112154 36090
rect 112154 36038 112156 36090
rect 112100 36036 112156 36038
rect 112204 36090 112260 36092
rect 112204 36038 112206 36090
rect 112206 36038 112258 36090
rect 112258 36038 112260 36090
rect 112204 36036 112260 36038
rect 111996 34522 112052 34524
rect 111996 34470 111998 34522
rect 111998 34470 112050 34522
rect 112050 34470 112052 34522
rect 111996 34468 112052 34470
rect 112100 34522 112156 34524
rect 112100 34470 112102 34522
rect 112102 34470 112154 34522
rect 112154 34470 112156 34522
rect 112100 34468 112156 34470
rect 112204 34522 112260 34524
rect 112204 34470 112206 34522
rect 112206 34470 112258 34522
rect 112258 34470 112260 34522
rect 112204 34468 112260 34470
rect 111996 32954 112052 32956
rect 111996 32902 111998 32954
rect 111998 32902 112050 32954
rect 112050 32902 112052 32954
rect 111996 32900 112052 32902
rect 112100 32954 112156 32956
rect 112100 32902 112102 32954
rect 112102 32902 112154 32954
rect 112154 32902 112156 32954
rect 112100 32900 112156 32902
rect 112204 32954 112260 32956
rect 112204 32902 112206 32954
rect 112206 32902 112258 32954
rect 112258 32902 112260 32954
rect 112204 32900 112260 32902
rect 111996 31386 112052 31388
rect 111996 31334 111998 31386
rect 111998 31334 112050 31386
rect 112050 31334 112052 31386
rect 111996 31332 112052 31334
rect 112100 31386 112156 31388
rect 112100 31334 112102 31386
rect 112102 31334 112154 31386
rect 112154 31334 112156 31386
rect 112100 31332 112156 31334
rect 112204 31386 112260 31388
rect 112204 31334 112206 31386
rect 112206 31334 112258 31386
rect 112258 31334 112260 31386
rect 112204 31332 112260 31334
rect 111996 29818 112052 29820
rect 111996 29766 111998 29818
rect 111998 29766 112050 29818
rect 112050 29766 112052 29818
rect 111996 29764 112052 29766
rect 112100 29818 112156 29820
rect 112100 29766 112102 29818
rect 112102 29766 112154 29818
rect 112154 29766 112156 29818
rect 112100 29764 112156 29766
rect 112204 29818 112260 29820
rect 112204 29766 112206 29818
rect 112206 29766 112258 29818
rect 112258 29766 112260 29818
rect 112204 29764 112260 29766
rect 111996 28250 112052 28252
rect 111996 28198 111998 28250
rect 111998 28198 112050 28250
rect 112050 28198 112052 28250
rect 111996 28196 112052 28198
rect 112100 28250 112156 28252
rect 112100 28198 112102 28250
rect 112102 28198 112154 28250
rect 112154 28198 112156 28250
rect 112100 28196 112156 28198
rect 112204 28250 112260 28252
rect 112204 28198 112206 28250
rect 112206 28198 112258 28250
rect 112258 28198 112260 28250
rect 112204 28196 112260 28198
rect 111996 26682 112052 26684
rect 111996 26630 111998 26682
rect 111998 26630 112050 26682
rect 112050 26630 112052 26682
rect 111996 26628 112052 26630
rect 112100 26682 112156 26684
rect 112100 26630 112102 26682
rect 112102 26630 112154 26682
rect 112154 26630 112156 26682
rect 112100 26628 112156 26630
rect 112204 26682 112260 26684
rect 112204 26630 112206 26682
rect 112206 26630 112258 26682
rect 112258 26630 112260 26682
rect 112204 26628 112260 26630
rect 111996 25114 112052 25116
rect 111996 25062 111998 25114
rect 111998 25062 112050 25114
rect 112050 25062 112052 25114
rect 111996 25060 112052 25062
rect 112100 25114 112156 25116
rect 112100 25062 112102 25114
rect 112102 25062 112154 25114
rect 112154 25062 112156 25114
rect 112100 25060 112156 25062
rect 112204 25114 112260 25116
rect 112204 25062 112206 25114
rect 112206 25062 112258 25114
rect 112258 25062 112260 25114
rect 112204 25060 112260 25062
rect 112364 23660 112420 23716
rect 111996 23546 112052 23548
rect 111996 23494 111998 23546
rect 111998 23494 112050 23546
rect 112050 23494 112052 23546
rect 111996 23492 112052 23494
rect 112100 23546 112156 23548
rect 112100 23494 112102 23546
rect 112102 23494 112154 23546
rect 112154 23494 112156 23546
rect 112100 23492 112156 23494
rect 112204 23546 112260 23548
rect 112204 23494 112206 23546
rect 112206 23494 112258 23546
rect 112258 23494 112260 23546
rect 112204 23492 112260 23494
rect 111996 21978 112052 21980
rect 111996 21926 111998 21978
rect 111998 21926 112050 21978
rect 112050 21926 112052 21978
rect 111996 21924 112052 21926
rect 112100 21978 112156 21980
rect 112100 21926 112102 21978
rect 112102 21926 112154 21978
rect 112154 21926 112156 21978
rect 112100 21924 112156 21926
rect 112204 21978 112260 21980
rect 112204 21926 112206 21978
rect 112206 21926 112258 21978
rect 112258 21926 112260 21978
rect 112204 21924 112260 21926
rect 111996 20410 112052 20412
rect 111996 20358 111998 20410
rect 111998 20358 112050 20410
rect 112050 20358 112052 20410
rect 111996 20356 112052 20358
rect 112100 20410 112156 20412
rect 112100 20358 112102 20410
rect 112102 20358 112154 20410
rect 112154 20358 112156 20410
rect 112100 20356 112156 20358
rect 112204 20410 112260 20412
rect 112204 20358 112206 20410
rect 112206 20358 112258 20410
rect 112258 20358 112260 20410
rect 112204 20356 112260 20358
rect 111996 18842 112052 18844
rect 111996 18790 111998 18842
rect 111998 18790 112050 18842
rect 112050 18790 112052 18842
rect 111996 18788 112052 18790
rect 112100 18842 112156 18844
rect 112100 18790 112102 18842
rect 112102 18790 112154 18842
rect 112154 18790 112156 18842
rect 112100 18788 112156 18790
rect 112204 18842 112260 18844
rect 112204 18790 112206 18842
rect 112206 18790 112258 18842
rect 112258 18790 112260 18842
rect 112204 18788 112260 18790
rect 111996 17274 112052 17276
rect 111996 17222 111998 17274
rect 111998 17222 112050 17274
rect 112050 17222 112052 17274
rect 111996 17220 112052 17222
rect 112100 17274 112156 17276
rect 112100 17222 112102 17274
rect 112102 17222 112154 17274
rect 112154 17222 112156 17274
rect 112100 17220 112156 17222
rect 112204 17274 112260 17276
rect 112204 17222 112206 17274
rect 112206 17222 112258 17274
rect 112258 17222 112260 17274
rect 112204 17220 112260 17222
rect 111996 15706 112052 15708
rect 111996 15654 111998 15706
rect 111998 15654 112050 15706
rect 112050 15654 112052 15706
rect 111996 15652 112052 15654
rect 112100 15706 112156 15708
rect 112100 15654 112102 15706
rect 112102 15654 112154 15706
rect 112154 15654 112156 15706
rect 112100 15652 112156 15654
rect 112204 15706 112260 15708
rect 112204 15654 112206 15706
rect 112206 15654 112258 15706
rect 112258 15654 112260 15706
rect 112204 15652 112260 15654
rect 111996 14138 112052 14140
rect 111996 14086 111998 14138
rect 111998 14086 112050 14138
rect 112050 14086 112052 14138
rect 111996 14084 112052 14086
rect 112100 14138 112156 14140
rect 112100 14086 112102 14138
rect 112102 14086 112154 14138
rect 112154 14086 112156 14138
rect 112100 14084 112156 14086
rect 112204 14138 112260 14140
rect 112204 14086 112206 14138
rect 112206 14086 112258 14138
rect 112258 14086 112260 14138
rect 112204 14084 112260 14086
rect 109228 13580 109284 13636
rect 111580 13580 111636 13636
rect 109452 12066 109508 12068
rect 109452 12014 109454 12066
rect 109454 12014 109506 12066
rect 109506 12014 109508 12066
rect 109452 12012 109508 12014
rect 111996 12570 112052 12572
rect 111996 12518 111998 12570
rect 111998 12518 112050 12570
rect 112050 12518 112052 12570
rect 111996 12516 112052 12518
rect 112100 12570 112156 12572
rect 112100 12518 112102 12570
rect 112102 12518 112154 12570
rect 112154 12518 112156 12570
rect 112100 12516 112156 12518
rect 112204 12570 112260 12572
rect 112204 12518 112206 12570
rect 112206 12518 112258 12570
rect 112258 12518 112260 12570
rect 112204 12516 112260 12518
rect 110796 11788 110852 11844
rect 109004 10556 109060 10612
rect 109900 11116 109956 11172
rect 110460 10780 110516 10836
rect 109900 10220 109956 10276
rect 110012 9548 110068 9604
rect 109116 9042 109172 9044
rect 109116 8990 109118 9042
rect 109118 8990 109170 9042
rect 109170 8990 109172 9042
rect 109116 8988 109172 8990
rect 110012 8988 110068 9044
rect 109900 8930 109956 8932
rect 109900 8878 109902 8930
rect 109902 8878 109954 8930
rect 109954 8878 109956 8930
rect 109900 8876 109956 8878
rect 109676 8652 109732 8708
rect 108780 8316 108836 8372
rect 109564 8540 109620 8596
rect 109340 8258 109396 8260
rect 109340 8206 109342 8258
rect 109342 8206 109394 8258
rect 109394 8206 109396 8258
rect 109340 8204 109396 8206
rect 109228 7980 109284 8036
rect 109004 7084 109060 7140
rect 108556 5292 108612 5348
rect 109452 7196 109508 7252
rect 109340 6466 109396 6468
rect 109340 6414 109342 6466
rect 109342 6414 109394 6466
rect 109394 6414 109396 6466
rect 109340 6412 109396 6414
rect 109564 6412 109620 6468
rect 109452 5740 109508 5796
rect 108892 4956 108948 5012
rect 108444 4172 108500 4228
rect 108444 3836 108500 3892
rect 109564 5068 109620 5124
rect 110012 8428 110068 8484
rect 110236 8764 110292 8820
rect 110236 7644 110292 7700
rect 110348 6524 110404 6580
rect 110348 5852 110404 5908
rect 110236 5122 110292 5124
rect 110236 5070 110238 5122
rect 110238 5070 110290 5122
rect 110290 5070 110292 5122
rect 110236 5068 110292 5070
rect 109900 4620 109956 4676
rect 109452 4060 109508 4116
rect 109564 4172 109620 4228
rect 109116 3612 109172 3668
rect 106876 3164 106932 3220
rect 107884 3388 107940 3444
rect 109004 3442 109060 3444
rect 109004 3390 109006 3442
rect 109006 3390 109058 3442
rect 109058 3390 109060 3442
rect 109004 3388 109060 3390
rect 110236 4226 110292 4228
rect 110236 4174 110238 4226
rect 110238 4174 110290 4226
rect 110290 4174 110292 4226
rect 110236 4172 110292 4174
rect 112140 12066 112196 12068
rect 112140 12014 112142 12066
rect 112142 12014 112194 12066
rect 112194 12014 112196 12066
rect 112140 12012 112196 12014
rect 111580 11788 111636 11844
rect 110796 8540 110852 8596
rect 111132 7980 111188 8036
rect 110796 7474 110852 7476
rect 110796 7422 110798 7474
rect 110798 7422 110850 7474
rect 110850 7422 110852 7474
rect 110796 7420 110852 7422
rect 111996 11002 112052 11004
rect 111996 10950 111998 11002
rect 111998 10950 112050 11002
rect 112050 10950 112052 11002
rect 111996 10948 112052 10950
rect 112100 11002 112156 11004
rect 112100 10950 112102 11002
rect 112102 10950 112154 11002
rect 112154 10950 112156 11002
rect 112100 10948 112156 10950
rect 112204 11002 112260 11004
rect 112204 10950 112206 11002
rect 112206 10950 112258 11002
rect 112258 10950 112260 11002
rect 112204 10948 112260 10950
rect 112028 10498 112084 10500
rect 112028 10446 112030 10498
rect 112030 10446 112082 10498
rect 112082 10446 112084 10498
rect 112028 10444 112084 10446
rect 112140 9996 112196 10052
rect 111692 7756 111748 7812
rect 111804 9884 111860 9940
rect 111580 7308 111636 7364
rect 111244 6972 111300 7028
rect 110572 4844 110628 4900
rect 110460 4620 110516 4676
rect 110796 6300 110852 6356
rect 110796 5852 110852 5908
rect 111020 5740 111076 5796
rect 111132 6412 111188 6468
rect 111132 5516 111188 5572
rect 111356 5404 111412 5460
rect 111356 4396 111412 4452
rect 111468 5346 111524 5348
rect 111468 5294 111470 5346
rect 111470 5294 111522 5346
rect 111522 5294 111524 5346
rect 111468 5292 111524 5294
rect 111468 4284 111524 4340
rect 112140 9660 112196 9716
rect 111996 9434 112052 9436
rect 111996 9382 111998 9434
rect 111998 9382 112050 9434
rect 112050 9382 112052 9434
rect 111996 9380 112052 9382
rect 112100 9434 112156 9436
rect 112100 9382 112102 9434
rect 112102 9382 112154 9434
rect 112154 9382 112156 9434
rect 112100 9380 112156 9382
rect 112204 9434 112260 9436
rect 112204 9382 112206 9434
rect 112206 9382 112258 9434
rect 112258 9382 112260 9434
rect 112204 9380 112260 9382
rect 112028 8988 112084 9044
rect 112252 8092 112308 8148
rect 111996 7866 112052 7868
rect 111996 7814 111998 7866
rect 111998 7814 112050 7866
rect 112050 7814 112052 7866
rect 111996 7812 112052 7814
rect 112100 7866 112156 7868
rect 112100 7814 112102 7866
rect 112102 7814 112154 7866
rect 112154 7814 112156 7866
rect 112100 7812 112156 7814
rect 112204 7866 112260 7868
rect 112204 7814 112206 7866
rect 112206 7814 112258 7866
rect 112258 7814 112260 7866
rect 112204 7812 112260 7814
rect 113596 19292 113652 19348
rect 113260 16828 113316 16884
rect 112588 11788 112644 11844
rect 113148 11170 113204 11172
rect 113148 11118 113150 11170
rect 113150 11118 113202 11170
rect 113202 11118 113204 11170
rect 113148 11116 113204 11118
rect 112700 11004 112756 11060
rect 113148 10220 113204 10276
rect 113596 10108 113652 10164
rect 112812 9602 112868 9604
rect 112812 9550 112814 9602
rect 112814 9550 112866 9602
rect 112866 9550 112868 9602
rect 112812 9548 112868 9550
rect 113036 9154 113092 9156
rect 113036 9102 113038 9154
rect 113038 9102 113090 9154
rect 113090 9102 113092 9154
rect 113036 9100 113092 9102
rect 113260 8370 113316 8372
rect 113260 8318 113262 8370
rect 113262 8318 113314 8370
rect 113314 8318 113316 8370
rect 113260 8316 113316 8318
rect 112588 7980 112644 8036
rect 112364 7756 112420 7812
rect 112812 7868 112868 7924
rect 112028 7308 112084 7364
rect 112812 7196 112868 7252
rect 112364 6972 112420 7028
rect 112140 6690 112196 6692
rect 112140 6638 112142 6690
rect 112142 6638 112194 6690
rect 112194 6638 112196 6690
rect 112140 6636 112196 6638
rect 111996 6298 112052 6300
rect 111996 6246 111998 6298
rect 111998 6246 112050 6298
rect 112050 6246 112052 6298
rect 111996 6244 112052 6246
rect 112100 6298 112156 6300
rect 112100 6246 112102 6298
rect 112102 6246 112154 6298
rect 112154 6246 112156 6298
rect 112100 6244 112156 6246
rect 112204 6298 112260 6300
rect 112204 6246 112206 6298
rect 112206 6246 112258 6298
rect 112258 6246 112260 6298
rect 112204 6244 112260 6246
rect 112588 5964 112644 6020
rect 112252 5292 112308 5348
rect 112700 5852 112756 5908
rect 111996 4730 112052 4732
rect 111996 4678 111998 4730
rect 111998 4678 112050 4730
rect 112050 4678 112052 4730
rect 111996 4676 112052 4678
rect 112100 4730 112156 4732
rect 112100 4678 112102 4730
rect 112102 4678 112154 4730
rect 112154 4678 112156 4730
rect 112100 4676 112156 4678
rect 112204 4730 112260 4732
rect 112204 4678 112206 4730
rect 112206 4678 112258 4730
rect 112258 4678 112260 4730
rect 112588 4732 112644 4788
rect 112204 4676 112260 4678
rect 110796 3724 110852 3780
rect 110796 2268 110852 2324
rect 111244 3388 111300 3444
rect 112364 3500 112420 3556
rect 111916 3442 111972 3444
rect 111916 3390 111918 3442
rect 111918 3390 111970 3442
rect 111970 3390 111972 3442
rect 111916 3388 111972 3390
rect 111996 3162 112052 3164
rect 111996 3110 111998 3162
rect 111998 3110 112050 3162
rect 112050 3110 112052 3162
rect 111996 3108 112052 3110
rect 112100 3162 112156 3164
rect 112100 3110 112102 3162
rect 112102 3110 112154 3162
rect 112154 3110 112156 3162
rect 112100 3108 112156 3110
rect 112204 3162 112260 3164
rect 112204 3110 112206 3162
rect 112206 3110 112258 3162
rect 112258 3110 112260 3162
rect 112204 3108 112260 3110
rect 113484 7308 113540 7364
rect 113036 6578 113092 6580
rect 113036 6526 113038 6578
rect 113038 6526 113090 6578
rect 113090 6526 113092 6578
rect 113036 6524 113092 6526
rect 113372 6188 113428 6244
rect 113148 5906 113204 5908
rect 113148 5854 113150 5906
rect 113150 5854 113202 5906
rect 113202 5854 113204 5906
rect 113148 5852 113204 5854
rect 113484 6076 113540 6132
rect 120540 116508 120596 116564
rect 121436 116562 121492 116564
rect 121436 116510 121438 116562
rect 121438 116510 121490 116562
rect 121490 116510 121492 116562
rect 121436 116508 121492 116510
rect 125244 116620 125300 116676
rect 126028 116620 126084 116676
rect 122108 116508 122164 116564
rect 124012 116562 124068 116564
rect 124012 116510 124014 116562
rect 124014 116510 124066 116562
rect 124066 116510 124068 116562
rect 124012 116508 124068 116510
rect 127356 116842 127412 116844
rect 127356 116790 127358 116842
rect 127358 116790 127410 116842
rect 127410 116790 127412 116842
rect 127356 116788 127412 116790
rect 127460 116842 127516 116844
rect 127460 116790 127462 116842
rect 127462 116790 127514 116842
rect 127514 116790 127516 116842
rect 127460 116788 127516 116790
rect 127564 116842 127620 116844
rect 127564 116790 127566 116842
rect 127566 116790 127618 116842
rect 127618 116790 127620 116842
rect 127564 116788 127620 116790
rect 126812 116508 126868 116564
rect 127932 116562 127988 116564
rect 127932 116510 127934 116562
rect 127934 116510 127986 116562
rect 127986 116510 127988 116562
rect 127932 116508 127988 116510
rect 129948 116508 130004 116564
rect 120092 116396 120148 116452
rect 118972 116172 119028 116228
rect 117404 115724 117460 115780
rect 118524 115778 118580 115780
rect 118524 115726 118526 115778
rect 118526 115726 118578 115778
rect 118578 115726 118580 115778
rect 118524 115724 118580 115726
rect 114940 115666 114996 115668
rect 114940 115614 114942 115666
rect 114942 115614 114994 115666
rect 114994 115614 114996 115666
rect 114940 115612 114996 115614
rect 115500 115666 115556 115668
rect 115500 115614 115502 115666
rect 115502 115614 115554 115666
rect 115554 115614 115556 115666
rect 115500 115612 115556 115614
rect 114380 115500 114436 115556
rect 115052 20748 115108 20804
rect 114828 19740 114884 19796
rect 113932 9772 113988 9828
rect 114156 17612 114212 17668
rect 114268 17052 114324 17108
rect 114716 12348 114772 12404
rect 114716 11170 114772 11172
rect 114716 11118 114718 11170
rect 114718 11118 114770 11170
rect 114770 11118 114772 11170
rect 114716 11116 114772 11118
rect 114268 10668 114324 10724
rect 114268 10108 114324 10164
rect 114156 9938 114212 9940
rect 114156 9886 114158 9938
rect 114158 9886 114210 9938
rect 114210 9886 114212 9938
rect 114156 9884 114212 9886
rect 114492 9660 114548 9716
rect 114380 9266 114436 9268
rect 114380 9214 114382 9266
rect 114382 9214 114434 9266
rect 114434 9214 114436 9266
rect 114380 9212 114436 9214
rect 113708 8652 113764 8708
rect 113708 8146 113764 8148
rect 113708 8094 113710 8146
rect 113710 8094 113762 8146
rect 113762 8094 113764 8146
rect 113708 8092 113764 8094
rect 113596 5794 113652 5796
rect 113596 5742 113598 5794
rect 113598 5742 113650 5794
rect 113650 5742 113652 5794
rect 113596 5740 113652 5742
rect 114044 8652 114100 8708
rect 113820 7308 113876 7364
rect 113932 7196 113988 7252
rect 118300 24108 118356 24164
rect 115836 19292 115892 19348
rect 115276 14364 115332 14420
rect 115276 11116 115332 11172
rect 115500 11788 115556 11844
rect 115164 9884 115220 9940
rect 114940 9212 114996 9268
rect 114716 8652 114772 8708
rect 114492 8428 114548 8484
rect 114156 8034 114212 8036
rect 114156 7982 114158 8034
rect 114158 7982 114210 8034
rect 114210 7982 114212 8034
rect 114156 7980 114212 7982
rect 114380 7698 114436 7700
rect 114380 7646 114382 7698
rect 114382 7646 114434 7698
rect 114434 7646 114436 7698
rect 114380 7644 114436 7646
rect 114268 7308 114324 7364
rect 114044 6636 114100 6692
rect 113708 5404 113764 5460
rect 114156 7196 114212 7252
rect 114044 6130 114100 6132
rect 114044 6078 114046 6130
rect 114046 6078 114098 6130
rect 114098 6078 114100 6130
rect 114044 6076 114100 6078
rect 113820 5516 113876 5572
rect 113036 5180 113092 5236
rect 113932 5404 113988 5460
rect 113372 4620 113428 4676
rect 113260 4562 113316 4564
rect 113260 4510 113262 4562
rect 113262 4510 113314 4562
rect 113314 4510 113316 4562
rect 113260 4508 113316 4510
rect 113708 4508 113764 4564
rect 113932 4844 113988 4900
rect 114716 8204 114772 8260
rect 114716 7644 114772 7700
rect 114828 7980 114884 8036
rect 114716 7420 114772 7476
rect 114268 6412 114324 6468
rect 114604 4396 114660 4452
rect 114492 4226 114548 4228
rect 114492 4174 114494 4226
rect 114494 4174 114546 4226
rect 114546 4174 114548 4226
rect 114492 4172 114548 4174
rect 112924 3612 112980 3668
rect 112700 2716 112756 2772
rect 111804 1372 111860 1428
rect 114044 3666 114100 3668
rect 114044 3614 114046 3666
rect 114046 3614 114098 3666
rect 114098 3614 114100 3666
rect 114044 3612 114100 3614
rect 113372 3554 113428 3556
rect 113372 3502 113374 3554
rect 113374 3502 113426 3554
rect 113426 3502 113428 3554
rect 113372 3500 113428 3502
rect 114492 1372 114548 1428
rect 114604 3388 114660 3444
rect 114828 6300 114884 6356
rect 115164 8204 115220 8260
rect 115164 7196 115220 7252
rect 115052 6188 115108 6244
rect 115164 6972 115220 7028
rect 114828 5068 114884 5124
rect 114940 5964 114996 6020
rect 114940 5292 114996 5348
rect 115612 10668 115668 10724
rect 115500 9324 115556 9380
rect 115500 8988 115556 9044
rect 116396 15820 116452 15876
rect 115948 10108 116004 10164
rect 116060 10332 116116 10388
rect 116396 9996 116452 10052
rect 115836 9212 115892 9268
rect 115948 9324 116004 9380
rect 115724 8316 115780 8372
rect 115836 8876 115892 8932
rect 115724 8034 115780 8036
rect 115724 7982 115726 8034
rect 115726 7982 115778 8034
rect 115778 7982 115780 8034
rect 115724 7980 115780 7982
rect 115388 7474 115444 7476
rect 115388 7422 115390 7474
rect 115390 7422 115442 7474
rect 115442 7422 115444 7474
rect 115388 7420 115444 7422
rect 115500 6972 115556 7028
rect 116396 9100 116452 9156
rect 116060 8258 116116 8260
rect 116060 8206 116062 8258
rect 116062 8206 116114 8258
rect 116114 8206 116116 8258
rect 116060 8204 116116 8206
rect 117180 12012 117236 12068
rect 116732 11116 116788 11172
rect 116620 9660 116676 9716
rect 117404 10780 117460 10836
rect 117292 10498 117348 10500
rect 117292 10446 117294 10498
rect 117294 10446 117346 10498
rect 117346 10446 117348 10498
rect 117292 10444 117348 10446
rect 116732 8652 116788 8708
rect 116508 8092 116564 8148
rect 116732 8092 116788 8148
rect 115948 7586 116004 7588
rect 115948 7534 115950 7586
rect 115950 7534 116002 7586
rect 116002 7534 116004 7586
rect 115948 7532 116004 7534
rect 115724 7420 115780 7476
rect 115836 7196 115892 7252
rect 115724 5068 115780 5124
rect 115612 4844 115668 4900
rect 115724 4620 115780 4676
rect 115164 4172 115220 4228
rect 115500 4172 115556 4228
rect 115948 6636 116004 6692
rect 116172 7868 116228 7924
rect 116284 6466 116340 6468
rect 116284 6414 116286 6466
rect 116286 6414 116338 6466
rect 116338 6414 116340 6466
rect 116284 6412 116340 6414
rect 116396 5964 116452 6020
rect 116620 6636 116676 6692
rect 116060 5292 116116 5348
rect 115948 4732 116004 4788
rect 116060 4508 116116 4564
rect 116172 4450 116228 4452
rect 116172 4398 116174 4450
rect 116174 4398 116226 4450
rect 116226 4398 116228 4450
rect 116172 4396 116228 4398
rect 117292 9714 117348 9716
rect 117292 9662 117294 9714
rect 117294 9662 117346 9714
rect 117346 9662 117348 9714
rect 117292 9660 117348 9662
rect 116956 8258 117012 8260
rect 116956 8206 116958 8258
rect 116958 8206 117010 8258
rect 117010 8206 117012 8258
rect 116956 8204 117012 8206
rect 117180 9154 117236 9156
rect 117180 9102 117182 9154
rect 117182 9102 117234 9154
rect 117234 9102 117236 9154
rect 117180 9100 117236 9102
rect 117516 9154 117572 9156
rect 117516 9102 117518 9154
rect 117518 9102 117570 9154
rect 117570 9102 117572 9154
rect 117516 9100 117572 9102
rect 117404 8652 117460 8708
rect 117292 8540 117348 8596
rect 116956 6300 117012 6356
rect 117180 8316 117236 8372
rect 117068 5292 117124 5348
rect 116956 4060 117012 4116
rect 116396 3836 116452 3892
rect 116284 3612 116340 3668
rect 114716 2156 114772 2212
rect 117292 7084 117348 7140
rect 117628 7420 117684 7476
rect 117404 6748 117460 6804
rect 118188 10498 118244 10500
rect 118188 10446 118190 10498
rect 118190 10446 118242 10498
rect 118242 10446 118244 10498
rect 118188 10444 118244 10446
rect 117964 8876 118020 8932
rect 117964 8428 118020 8484
rect 118188 10220 118244 10276
rect 118076 8092 118132 8148
rect 118412 9660 118468 9716
rect 118300 8034 118356 8036
rect 118300 7982 118302 8034
rect 118302 7982 118354 8034
rect 118354 7982 118356 8034
rect 118300 7980 118356 7982
rect 117852 6748 117908 6804
rect 118188 7196 118244 7252
rect 117628 6018 117684 6020
rect 117628 5966 117630 6018
rect 117630 5966 117682 6018
rect 117682 5966 117684 6018
rect 117628 5964 117684 5966
rect 117740 5682 117796 5684
rect 117740 5630 117742 5682
rect 117742 5630 117794 5682
rect 117794 5630 117796 5682
rect 117740 5628 117796 5630
rect 117516 5292 117572 5348
rect 117404 5068 117460 5124
rect 117516 4844 117572 4900
rect 117404 4562 117460 4564
rect 117404 4510 117406 4562
rect 117406 4510 117458 4562
rect 117458 4510 117460 4562
rect 117404 4508 117460 4510
rect 117628 4732 117684 4788
rect 118076 5852 118132 5908
rect 117964 4284 118020 4340
rect 117964 3666 118020 3668
rect 117964 3614 117966 3666
rect 117966 3614 118018 3666
rect 118018 3614 118020 3666
rect 117964 3612 118020 3614
rect 116396 3442 116452 3444
rect 116396 3390 116398 3442
rect 116398 3390 116450 3442
rect 116450 3390 116452 3442
rect 116396 3388 116452 3390
rect 117964 3388 118020 3444
rect 118412 7756 118468 7812
rect 118636 9548 118692 9604
rect 118748 8316 118804 8372
rect 118524 7644 118580 7700
rect 118748 7980 118804 8036
rect 118524 7420 118580 7476
rect 118860 7868 118916 7924
rect 118860 7532 118916 7588
rect 118748 7474 118804 7476
rect 118748 7422 118750 7474
rect 118750 7422 118802 7474
rect 118802 7422 118804 7474
rect 118748 7420 118804 7422
rect 122556 116226 122612 116228
rect 122556 116174 122558 116226
rect 122558 116174 122610 116226
rect 122610 116174 122612 116226
rect 122556 116172 122612 116174
rect 123340 116172 123396 116228
rect 129836 116396 129892 116452
rect 120316 115666 120372 115668
rect 120316 115614 120318 115666
rect 120318 115614 120370 115666
rect 120370 115614 120372 115666
rect 120316 115612 120372 115614
rect 121324 115666 121380 115668
rect 121324 115614 121326 115666
rect 121326 115614 121378 115666
rect 121378 115614 121380 115666
rect 121324 115612 121380 115614
rect 124236 115666 124292 115668
rect 124236 115614 124238 115666
rect 124238 115614 124290 115666
rect 124290 115614 124292 115666
rect 124236 115612 124292 115614
rect 124796 115666 124852 115668
rect 124796 115614 124798 115666
rect 124798 115614 124850 115666
rect 124850 115614 124852 115666
rect 124796 115612 124852 115614
rect 125244 115500 125300 115556
rect 120540 27020 120596 27076
rect 120764 26908 120820 26964
rect 124572 23996 124628 24052
rect 123340 22204 123396 22260
rect 120092 11788 120148 11844
rect 119308 11116 119364 11172
rect 119084 11004 119140 11060
rect 120204 10668 120260 10724
rect 119308 9996 119364 10052
rect 119980 10332 120036 10388
rect 119196 9714 119252 9716
rect 119196 9662 119198 9714
rect 119198 9662 119250 9714
rect 119250 9662 119252 9714
rect 119196 9660 119252 9662
rect 119308 9100 119364 9156
rect 119196 8930 119252 8932
rect 119196 8878 119198 8930
rect 119198 8878 119250 8930
rect 119250 8878 119252 8930
rect 119196 8876 119252 8878
rect 119084 8204 119140 8260
rect 119196 8652 119252 8708
rect 118972 7308 119028 7364
rect 118972 7084 119028 7140
rect 118748 6466 118804 6468
rect 118748 6414 118750 6466
rect 118750 6414 118802 6466
rect 118802 6414 118804 6466
rect 118748 6412 118804 6414
rect 118636 5852 118692 5908
rect 118748 5682 118804 5684
rect 118748 5630 118750 5682
rect 118750 5630 118802 5682
rect 118802 5630 118804 5682
rect 118748 5628 118804 5630
rect 118524 5068 118580 5124
rect 118636 5516 118692 5572
rect 119084 6802 119140 6804
rect 119084 6750 119086 6802
rect 119086 6750 119138 6802
rect 119138 6750 119140 6802
rect 119084 6748 119140 6750
rect 118972 5068 119028 5124
rect 119084 5516 119140 5572
rect 118860 4284 118916 4340
rect 118636 4226 118692 4228
rect 118636 4174 118638 4226
rect 118638 4174 118690 4226
rect 118690 4174 118692 4226
rect 118636 4172 118692 4174
rect 118076 3276 118132 3332
rect 119868 8652 119924 8708
rect 120204 10332 120260 10388
rect 120316 9212 120372 9268
rect 119980 8316 120036 8372
rect 119644 8258 119700 8260
rect 119644 8206 119646 8258
rect 119646 8206 119698 8258
rect 119698 8206 119700 8258
rect 119644 8204 119700 8206
rect 119756 7980 119812 8036
rect 119532 7756 119588 7812
rect 119420 7362 119476 7364
rect 119420 7310 119422 7362
rect 119422 7310 119474 7362
rect 119474 7310 119476 7362
rect 119420 7308 119476 7310
rect 119308 6860 119364 6916
rect 119644 7532 119700 7588
rect 119532 6972 119588 7028
rect 119868 6860 119924 6916
rect 119756 6748 119812 6804
rect 119868 6300 119924 6356
rect 119868 5906 119924 5908
rect 119868 5854 119870 5906
rect 119870 5854 119922 5906
rect 119922 5854 119924 5906
rect 119868 5852 119924 5854
rect 119532 5682 119588 5684
rect 119532 5630 119534 5682
rect 119534 5630 119586 5682
rect 119586 5630 119588 5682
rect 119532 5628 119588 5630
rect 119868 5234 119924 5236
rect 119868 5182 119870 5234
rect 119870 5182 119922 5234
rect 119922 5182 119924 5234
rect 119868 5180 119924 5182
rect 120092 6860 120148 6916
rect 123228 17500 123284 17556
rect 120876 9212 120932 9268
rect 121884 9266 121940 9268
rect 121884 9214 121886 9266
rect 121886 9214 121938 9266
rect 121938 9214 121940 9266
rect 121884 9212 121940 9214
rect 120988 8988 121044 9044
rect 121548 9042 121604 9044
rect 121548 8990 121550 9042
rect 121550 8990 121602 9042
rect 121602 8990 121604 9042
rect 121548 8988 121604 8990
rect 120428 7980 120484 8036
rect 120316 7362 120372 7364
rect 120316 7310 120318 7362
rect 120318 7310 120370 7362
rect 120370 7310 120372 7362
rect 120316 7308 120372 7310
rect 120204 6802 120260 6804
rect 120204 6750 120206 6802
rect 120206 6750 120258 6802
rect 120258 6750 120260 6802
rect 120204 6748 120260 6750
rect 120092 6412 120148 6468
rect 119756 5068 119812 5124
rect 119420 4844 119476 4900
rect 119420 4450 119476 4452
rect 119420 4398 119422 4450
rect 119422 4398 119474 4450
rect 119474 4398 119476 4450
rect 119420 4396 119476 4398
rect 120428 6300 120484 6356
rect 120204 4396 120260 4452
rect 120988 8316 121044 8372
rect 120652 8258 120708 8260
rect 120652 8206 120654 8258
rect 120654 8206 120706 8258
rect 120706 8206 120708 8258
rect 120652 8204 120708 8206
rect 120764 7980 120820 8036
rect 120652 6636 120708 6692
rect 120652 6300 120708 6356
rect 121212 8092 121268 8148
rect 121100 7084 121156 7140
rect 121436 7586 121492 7588
rect 121436 7534 121438 7586
rect 121438 7534 121490 7586
rect 121490 7534 121492 7586
rect 121436 7532 121492 7534
rect 120876 5068 120932 5124
rect 121324 7308 121380 7364
rect 120876 4508 120932 4564
rect 119868 4338 119924 4340
rect 119868 4286 119870 4338
rect 119870 4286 119922 4338
rect 119922 4286 119924 4338
rect 119868 4284 119924 4286
rect 119644 3836 119700 3892
rect 119196 2828 119252 2884
rect 119644 3276 119700 3332
rect 120092 3052 120148 3108
rect 120204 3724 120260 3780
rect 120764 3612 120820 3668
rect 120316 3442 120372 3444
rect 120316 3390 120318 3442
rect 120318 3390 120370 3442
rect 120370 3390 120372 3442
rect 120316 3388 120372 3390
rect 121100 5794 121156 5796
rect 121100 5742 121102 5794
rect 121102 5742 121154 5794
rect 121154 5742 121156 5794
rect 121100 5740 121156 5742
rect 121100 4844 121156 4900
rect 121436 5794 121492 5796
rect 121436 5742 121438 5794
rect 121438 5742 121490 5794
rect 121490 5742 121492 5794
rect 121436 5740 121492 5742
rect 121212 4620 121268 4676
rect 121436 4620 121492 4676
rect 121324 4562 121380 4564
rect 121324 4510 121326 4562
rect 121326 4510 121378 4562
rect 121378 4510 121380 4562
rect 121324 4508 121380 4510
rect 121212 4338 121268 4340
rect 121212 4286 121214 4338
rect 121214 4286 121266 4338
rect 121266 4286 121268 4338
rect 121212 4284 121268 4286
rect 121996 8034 122052 8036
rect 121996 7982 121998 8034
rect 121998 7982 122050 8034
rect 122050 7982 122052 8034
rect 121996 7980 122052 7982
rect 121884 7868 121940 7924
rect 121660 5516 121716 5572
rect 121772 6972 121828 7028
rect 121660 5292 121716 5348
rect 122220 7756 122276 7812
rect 121996 7362 122052 7364
rect 121996 7310 121998 7362
rect 121998 7310 122050 7362
rect 122050 7310 122052 7362
rect 121996 7308 122052 7310
rect 121996 6860 122052 6916
rect 121996 6466 122052 6468
rect 121996 6414 121998 6466
rect 121998 6414 122050 6466
rect 122050 6414 122052 6466
rect 121996 6412 122052 6414
rect 121996 5964 122052 6020
rect 121996 5794 122052 5796
rect 121996 5742 121998 5794
rect 121998 5742 122050 5794
rect 122050 5742 122052 5794
rect 121996 5740 122052 5742
rect 121884 5234 121940 5236
rect 121884 5182 121886 5234
rect 121886 5182 121938 5234
rect 121938 5182 121940 5234
rect 121884 5180 121940 5182
rect 121772 4956 121828 5012
rect 121548 4396 121604 4452
rect 121660 4508 121716 4564
rect 121548 4060 121604 4116
rect 121436 3836 121492 3892
rect 121212 3554 121268 3556
rect 121212 3502 121214 3554
rect 121214 3502 121266 3554
rect 121266 3502 121268 3554
rect 121212 3500 121268 3502
rect 120988 3388 121044 3444
rect 122108 5404 122164 5460
rect 122108 4956 122164 5012
rect 123228 7698 123284 7700
rect 123228 7646 123230 7698
rect 123230 7646 123282 7698
rect 123282 7646 123284 7698
rect 123228 7644 123284 7646
rect 122444 7420 122500 7476
rect 122444 7196 122500 7252
rect 122444 6690 122500 6692
rect 122444 6638 122446 6690
rect 122446 6638 122498 6690
rect 122498 6638 122500 6690
rect 122444 6636 122500 6638
rect 122332 6076 122388 6132
rect 122780 6636 122836 6692
rect 123452 8876 123508 8932
rect 124124 8764 124180 8820
rect 122668 5852 122724 5908
rect 122668 5292 122724 5348
rect 122780 6412 122836 6468
rect 122332 4338 122388 4340
rect 122332 4286 122334 4338
rect 122334 4286 122386 4338
rect 122386 4286 122388 4338
rect 122332 4284 122388 4286
rect 122220 4172 122276 4228
rect 121884 3612 121940 3668
rect 121772 3442 121828 3444
rect 121772 3390 121774 3442
rect 121774 3390 121826 3442
rect 121826 3390 121828 3442
rect 121772 3388 121828 3390
rect 122444 3330 122500 3332
rect 122444 3278 122446 3330
rect 122446 3278 122498 3330
rect 122498 3278 122500 3330
rect 122444 3276 122500 3278
rect 123900 8428 123956 8484
rect 123452 6748 123508 6804
rect 122892 5516 122948 5572
rect 122892 5068 122948 5124
rect 122668 4060 122724 4116
rect 122556 3164 122612 3220
rect 123340 6076 123396 6132
rect 123452 5346 123508 5348
rect 123452 5294 123454 5346
rect 123454 5294 123506 5346
rect 123506 5294 123508 5346
rect 123452 5292 123508 5294
rect 123228 3948 123284 4004
rect 123340 4844 123396 4900
rect 123900 6412 123956 6468
rect 123788 6188 123844 6244
rect 123788 6018 123844 6020
rect 123788 5966 123790 6018
rect 123790 5966 123842 6018
rect 123842 5966 123844 6018
rect 123788 5964 123844 5966
rect 123788 5628 123844 5684
rect 123676 5122 123732 5124
rect 123676 5070 123678 5122
rect 123678 5070 123730 5122
rect 123730 5070 123732 5122
rect 123676 5068 123732 5070
rect 123564 4620 123620 4676
rect 124236 8652 124292 8708
rect 124236 8092 124292 8148
rect 124236 6300 124292 6356
rect 123900 4620 123956 4676
rect 123564 4060 123620 4116
rect 124236 4956 124292 5012
rect 124124 4060 124180 4116
rect 123676 3836 123732 3892
rect 124124 3836 124180 3892
rect 123564 3388 123620 3444
rect 123228 1260 123284 1316
rect 124460 5292 124516 5348
rect 131180 116450 131236 116452
rect 131180 116398 131182 116450
rect 131182 116398 131234 116450
rect 131234 116398 131236 116450
rect 131180 116396 131236 116398
rect 131852 116562 131908 116564
rect 131852 116510 131854 116562
rect 131854 116510 131906 116562
rect 131906 116510 131908 116562
rect 131852 116508 131908 116510
rect 139356 116620 139412 116676
rect 140252 116620 140308 116676
rect 131516 115724 131572 115780
rect 132636 115778 132692 115780
rect 132636 115726 132638 115778
rect 132638 115726 132690 115778
rect 132690 115726 132692 115778
rect 132636 115724 132692 115726
rect 128940 115666 128996 115668
rect 128940 115614 128942 115666
rect 128942 115614 128994 115666
rect 128994 115614 128996 115666
rect 128940 115612 128996 115614
rect 129612 115666 129668 115668
rect 129612 115614 129614 115666
rect 129614 115614 129666 115666
rect 129666 115614 129668 115666
rect 129612 115612 129668 115614
rect 126924 115500 126980 115556
rect 133756 115666 133812 115668
rect 133756 115614 133758 115666
rect 133758 115614 133810 115666
rect 133810 115614 133812 115666
rect 133756 115612 133812 115614
rect 134316 115666 134372 115668
rect 134316 115614 134318 115666
rect 134318 115614 134370 115666
rect 134370 115614 134372 115666
rect 134316 115612 134372 115614
rect 127356 115274 127412 115276
rect 127356 115222 127358 115274
rect 127358 115222 127410 115274
rect 127410 115222 127412 115274
rect 127356 115220 127412 115222
rect 127460 115274 127516 115276
rect 127460 115222 127462 115274
rect 127462 115222 127514 115274
rect 127514 115222 127516 115274
rect 127460 115220 127516 115222
rect 127564 115274 127620 115276
rect 127564 115222 127566 115274
rect 127566 115222 127618 115274
rect 127618 115222 127620 115274
rect 127564 115220 127620 115222
rect 127356 113706 127412 113708
rect 127356 113654 127358 113706
rect 127358 113654 127410 113706
rect 127410 113654 127412 113706
rect 127356 113652 127412 113654
rect 127460 113706 127516 113708
rect 127460 113654 127462 113706
rect 127462 113654 127514 113706
rect 127514 113654 127516 113706
rect 127460 113652 127516 113654
rect 127564 113706 127620 113708
rect 127564 113654 127566 113706
rect 127566 113654 127618 113706
rect 127618 113654 127620 113706
rect 127564 113652 127620 113654
rect 127356 112138 127412 112140
rect 127356 112086 127358 112138
rect 127358 112086 127410 112138
rect 127410 112086 127412 112138
rect 127356 112084 127412 112086
rect 127460 112138 127516 112140
rect 127460 112086 127462 112138
rect 127462 112086 127514 112138
rect 127514 112086 127516 112138
rect 127460 112084 127516 112086
rect 127564 112138 127620 112140
rect 127564 112086 127566 112138
rect 127566 112086 127618 112138
rect 127618 112086 127620 112138
rect 127564 112084 127620 112086
rect 127356 110570 127412 110572
rect 127356 110518 127358 110570
rect 127358 110518 127410 110570
rect 127410 110518 127412 110570
rect 127356 110516 127412 110518
rect 127460 110570 127516 110572
rect 127460 110518 127462 110570
rect 127462 110518 127514 110570
rect 127514 110518 127516 110570
rect 127460 110516 127516 110518
rect 127564 110570 127620 110572
rect 127564 110518 127566 110570
rect 127566 110518 127618 110570
rect 127618 110518 127620 110570
rect 127564 110516 127620 110518
rect 127356 109002 127412 109004
rect 127356 108950 127358 109002
rect 127358 108950 127410 109002
rect 127410 108950 127412 109002
rect 127356 108948 127412 108950
rect 127460 109002 127516 109004
rect 127460 108950 127462 109002
rect 127462 108950 127514 109002
rect 127514 108950 127516 109002
rect 127460 108948 127516 108950
rect 127564 109002 127620 109004
rect 127564 108950 127566 109002
rect 127566 108950 127618 109002
rect 127618 108950 127620 109002
rect 127564 108948 127620 108950
rect 127356 107434 127412 107436
rect 127356 107382 127358 107434
rect 127358 107382 127410 107434
rect 127410 107382 127412 107434
rect 127356 107380 127412 107382
rect 127460 107434 127516 107436
rect 127460 107382 127462 107434
rect 127462 107382 127514 107434
rect 127514 107382 127516 107434
rect 127460 107380 127516 107382
rect 127564 107434 127620 107436
rect 127564 107382 127566 107434
rect 127566 107382 127618 107434
rect 127618 107382 127620 107434
rect 127564 107380 127620 107382
rect 127356 105866 127412 105868
rect 127356 105814 127358 105866
rect 127358 105814 127410 105866
rect 127410 105814 127412 105866
rect 127356 105812 127412 105814
rect 127460 105866 127516 105868
rect 127460 105814 127462 105866
rect 127462 105814 127514 105866
rect 127514 105814 127516 105866
rect 127460 105812 127516 105814
rect 127564 105866 127620 105868
rect 127564 105814 127566 105866
rect 127566 105814 127618 105866
rect 127618 105814 127620 105866
rect 127564 105812 127620 105814
rect 127356 104298 127412 104300
rect 127356 104246 127358 104298
rect 127358 104246 127410 104298
rect 127410 104246 127412 104298
rect 127356 104244 127412 104246
rect 127460 104298 127516 104300
rect 127460 104246 127462 104298
rect 127462 104246 127514 104298
rect 127514 104246 127516 104298
rect 127460 104244 127516 104246
rect 127564 104298 127620 104300
rect 127564 104246 127566 104298
rect 127566 104246 127618 104298
rect 127618 104246 127620 104298
rect 127564 104244 127620 104246
rect 127356 102730 127412 102732
rect 127356 102678 127358 102730
rect 127358 102678 127410 102730
rect 127410 102678 127412 102730
rect 127356 102676 127412 102678
rect 127460 102730 127516 102732
rect 127460 102678 127462 102730
rect 127462 102678 127514 102730
rect 127514 102678 127516 102730
rect 127460 102676 127516 102678
rect 127564 102730 127620 102732
rect 127564 102678 127566 102730
rect 127566 102678 127618 102730
rect 127618 102678 127620 102730
rect 127564 102676 127620 102678
rect 127356 101162 127412 101164
rect 127356 101110 127358 101162
rect 127358 101110 127410 101162
rect 127410 101110 127412 101162
rect 127356 101108 127412 101110
rect 127460 101162 127516 101164
rect 127460 101110 127462 101162
rect 127462 101110 127514 101162
rect 127514 101110 127516 101162
rect 127460 101108 127516 101110
rect 127564 101162 127620 101164
rect 127564 101110 127566 101162
rect 127566 101110 127618 101162
rect 127618 101110 127620 101162
rect 127564 101108 127620 101110
rect 127356 99594 127412 99596
rect 127356 99542 127358 99594
rect 127358 99542 127410 99594
rect 127410 99542 127412 99594
rect 127356 99540 127412 99542
rect 127460 99594 127516 99596
rect 127460 99542 127462 99594
rect 127462 99542 127514 99594
rect 127514 99542 127516 99594
rect 127460 99540 127516 99542
rect 127564 99594 127620 99596
rect 127564 99542 127566 99594
rect 127566 99542 127618 99594
rect 127618 99542 127620 99594
rect 127564 99540 127620 99542
rect 127356 98026 127412 98028
rect 127356 97974 127358 98026
rect 127358 97974 127410 98026
rect 127410 97974 127412 98026
rect 127356 97972 127412 97974
rect 127460 98026 127516 98028
rect 127460 97974 127462 98026
rect 127462 97974 127514 98026
rect 127514 97974 127516 98026
rect 127460 97972 127516 97974
rect 127564 98026 127620 98028
rect 127564 97974 127566 98026
rect 127566 97974 127618 98026
rect 127618 97974 127620 98026
rect 127564 97972 127620 97974
rect 127356 96458 127412 96460
rect 127356 96406 127358 96458
rect 127358 96406 127410 96458
rect 127410 96406 127412 96458
rect 127356 96404 127412 96406
rect 127460 96458 127516 96460
rect 127460 96406 127462 96458
rect 127462 96406 127514 96458
rect 127514 96406 127516 96458
rect 127460 96404 127516 96406
rect 127564 96458 127620 96460
rect 127564 96406 127566 96458
rect 127566 96406 127618 96458
rect 127618 96406 127620 96458
rect 127564 96404 127620 96406
rect 127356 94890 127412 94892
rect 127356 94838 127358 94890
rect 127358 94838 127410 94890
rect 127410 94838 127412 94890
rect 127356 94836 127412 94838
rect 127460 94890 127516 94892
rect 127460 94838 127462 94890
rect 127462 94838 127514 94890
rect 127514 94838 127516 94890
rect 127460 94836 127516 94838
rect 127564 94890 127620 94892
rect 127564 94838 127566 94890
rect 127566 94838 127618 94890
rect 127618 94838 127620 94890
rect 127564 94836 127620 94838
rect 127356 93322 127412 93324
rect 127356 93270 127358 93322
rect 127358 93270 127410 93322
rect 127410 93270 127412 93322
rect 127356 93268 127412 93270
rect 127460 93322 127516 93324
rect 127460 93270 127462 93322
rect 127462 93270 127514 93322
rect 127514 93270 127516 93322
rect 127460 93268 127516 93270
rect 127564 93322 127620 93324
rect 127564 93270 127566 93322
rect 127566 93270 127618 93322
rect 127618 93270 127620 93322
rect 127564 93268 127620 93270
rect 127356 91754 127412 91756
rect 127356 91702 127358 91754
rect 127358 91702 127410 91754
rect 127410 91702 127412 91754
rect 127356 91700 127412 91702
rect 127460 91754 127516 91756
rect 127460 91702 127462 91754
rect 127462 91702 127514 91754
rect 127514 91702 127516 91754
rect 127460 91700 127516 91702
rect 127564 91754 127620 91756
rect 127564 91702 127566 91754
rect 127566 91702 127618 91754
rect 127618 91702 127620 91754
rect 127564 91700 127620 91702
rect 127356 90186 127412 90188
rect 127356 90134 127358 90186
rect 127358 90134 127410 90186
rect 127410 90134 127412 90186
rect 127356 90132 127412 90134
rect 127460 90186 127516 90188
rect 127460 90134 127462 90186
rect 127462 90134 127514 90186
rect 127514 90134 127516 90186
rect 127460 90132 127516 90134
rect 127564 90186 127620 90188
rect 127564 90134 127566 90186
rect 127566 90134 127618 90186
rect 127618 90134 127620 90186
rect 127564 90132 127620 90134
rect 127356 88618 127412 88620
rect 127356 88566 127358 88618
rect 127358 88566 127410 88618
rect 127410 88566 127412 88618
rect 127356 88564 127412 88566
rect 127460 88618 127516 88620
rect 127460 88566 127462 88618
rect 127462 88566 127514 88618
rect 127514 88566 127516 88618
rect 127460 88564 127516 88566
rect 127564 88618 127620 88620
rect 127564 88566 127566 88618
rect 127566 88566 127618 88618
rect 127618 88566 127620 88618
rect 127564 88564 127620 88566
rect 127356 87050 127412 87052
rect 127356 86998 127358 87050
rect 127358 86998 127410 87050
rect 127410 86998 127412 87050
rect 127356 86996 127412 86998
rect 127460 87050 127516 87052
rect 127460 86998 127462 87050
rect 127462 86998 127514 87050
rect 127514 86998 127516 87050
rect 127460 86996 127516 86998
rect 127564 87050 127620 87052
rect 127564 86998 127566 87050
rect 127566 86998 127618 87050
rect 127618 86998 127620 87050
rect 127564 86996 127620 86998
rect 127356 85482 127412 85484
rect 127356 85430 127358 85482
rect 127358 85430 127410 85482
rect 127410 85430 127412 85482
rect 127356 85428 127412 85430
rect 127460 85482 127516 85484
rect 127460 85430 127462 85482
rect 127462 85430 127514 85482
rect 127514 85430 127516 85482
rect 127460 85428 127516 85430
rect 127564 85482 127620 85484
rect 127564 85430 127566 85482
rect 127566 85430 127618 85482
rect 127618 85430 127620 85482
rect 127564 85428 127620 85430
rect 127356 83914 127412 83916
rect 127356 83862 127358 83914
rect 127358 83862 127410 83914
rect 127410 83862 127412 83914
rect 127356 83860 127412 83862
rect 127460 83914 127516 83916
rect 127460 83862 127462 83914
rect 127462 83862 127514 83914
rect 127514 83862 127516 83914
rect 127460 83860 127516 83862
rect 127564 83914 127620 83916
rect 127564 83862 127566 83914
rect 127566 83862 127618 83914
rect 127618 83862 127620 83914
rect 127564 83860 127620 83862
rect 127356 82346 127412 82348
rect 127356 82294 127358 82346
rect 127358 82294 127410 82346
rect 127410 82294 127412 82346
rect 127356 82292 127412 82294
rect 127460 82346 127516 82348
rect 127460 82294 127462 82346
rect 127462 82294 127514 82346
rect 127514 82294 127516 82346
rect 127460 82292 127516 82294
rect 127564 82346 127620 82348
rect 127564 82294 127566 82346
rect 127566 82294 127618 82346
rect 127618 82294 127620 82346
rect 127564 82292 127620 82294
rect 127356 80778 127412 80780
rect 127356 80726 127358 80778
rect 127358 80726 127410 80778
rect 127410 80726 127412 80778
rect 127356 80724 127412 80726
rect 127460 80778 127516 80780
rect 127460 80726 127462 80778
rect 127462 80726 127514 80778
rect 127514 80726 127516 80778
rect 127460 80724 127516 80726
rect 127564 80778 127620 80780
rect 127564 80726 127566 80778
rect 127566 80726 127618 80778
rect 127618 80726 127620 80778
rect 127564 80724 127620 80726
rect 127356 79210 127412 79212
rect 127356 79158 127358 79210
rect 127358 79158 127410 79210
rect 127410 79158 127412 79210
rect 127356 79156 127412 79158
rect 127460 79210 127516 79212
rect 127460 79158 127462 79210
rect 127462 79158 127514 79210
rect 127514 79158 127516 79210
rect 127460 79156 127516 79158
rect 127564 79210 127620 79212
rect 127564 79158 127566 79210
rect 127566 79158 127618 79210
rect 127618 79158 127620 79210
rect 127564 79156 127620 79158
rect 127356 77642 127412 77644
rect 127356 77590 127358 77642
rect 127358 77590 127410 77642
rect 127410 77590 127412 77642
rect 127356 77588 127412 77590
rect 127460 77642 127516 77644
rect 127460 77590 127462 77642
rect 127462 77590 127514 77642
rect 127514 77590 127516 77642
rect 127460 77588 127516 77590
rect 127564 77642 127620 77644
rect 127564 77590 127566 77642
rect 127566 77590 127618 77642
rect 127618 77590 127620 77642
rect 127564 77588 127620 77590
rect 127356 76074 127412 76076
rect 127356 76022 127358 76074
rect 127358 76022 127410 76074
rect 127410 76022 127412 76074
rect 127356 76020 127412 76022
rect 127460 76074 127516 76076
rect 127460 76022 127462 76074
rect 127462 76022 127514 76074
rect 127514 76022 127516 76074
rect 127460 76020 127516 76022
rect 127564 76074 127620 76076
rect 127564 76022 127566 76074
rect 127566 76022 127618 76074
rect 127618 76022 127620 76074
rect 127564 76020 127620 76022
rect 127356 74506 127412 74508
rect 127356 74454 127358 74506
rect 127358 74454 127410 74506
rect 127410 74454 127412 74506
rect 127356 74452 127412 74454
rect 127460 74506 127516 74508
rect 127460 74454 127462 74506
rect 127462 74454 127514 74506
rect 127514 74454 127516 74506
rect 127460 74452 127516 74454
rect 127564 74506 127620 74508
rect 127564 74454 127566 74506
rect 127566 74454 127618 74506
rect 127618 74454 127620 74506
rect 127564 74452 127620 74454
rect 127356 72938 127412 72940
rect 127356 72886 127358 72938
rect 127358 72886 127410 72938
rect 127410 72886 127412 72938
rect 127356 72884 127412 72886
rect 127460 72938 127516 72940
rect 127460 72886 127462 72938
rect 127462 72886 127514 72938
rect 127514 72886 127516 72938
rect 127460 72884 127516 72886
rect 127564 72938 127620 72940
rect 127564 72886 127566 72938
rect 127566 72886 127618 72938
rect 127618 72886 127620 72938
rect 127564 72884 127620 72886
rect 127356 71370 127412 71372
rect 127356 71318 127358 71370
rect 127358 71318 127410 71370
rect 127410 71318 127412 71370
rect 127356 71316 127412 71318
rect 127460 71370 127516 71372
rect 127460 71318 127462 71370
rect 127462 71318 127514 71370
rect 127514 71318 127516 71370
rect 127460 71316 127516 71318
rect 127564 71370 127620 71372
rect 127564 71318 127566 71370
rect 127566 71318 127618 71370
rect 127618 71318 127620 71370
rect 127564 71316 127620 71318
rect 127356 69802 127412 69804
rect 127356 69750 127358 69802
rect 127358 69750 127410 69802
rect 127410 69750 127412 69802
rect 127356 69748 127412 69750
rect 127460 69802 127516 69804
rect 127460 69750 127462 69802
rect 127462 69750 127514 69802
rect 127514 69750 127516 69802
rect 127460 69748 127516 69750
rect 127564 69802 127620 69804
rect 127564 69750 127566 69802
rect 127566 69750 127618 69802
rect 127618 69750 127620 69802
rect 127564 69748 127620 69750
rect 127356 68234 127412 68236
rect 127356 68182 127358 68234
rect 127358 68182 127410 68234
rect 127410 68182 127412 68234
rect 127356 68180 127412 68182
rect 127460 68234 127516 68236
rect 127460 68182 127462 68234
rect 127462 68182 127514 68234
rect 127514 68182 127516 68234
rect 127460 68180 127516 68182
rect 127564 68234 127620 68236
rect 127564 68182 127566 68234
rect 127566 68182 127618 68234
rect 127618 68182 127620 68234
rect 127564 68180 127620 68182
rect 127356 66666 127412 66668
rect 127356 66614 127358 66666
rect 127358 66614 127410 66666
rect 127410 66614 127412 66666
rect 127356 66612 127412 66614
rect 127460 66666 127516 66668
rect 127460 66614 127462 66666
rect 127462 66614 127514 66666
rect 127514 66614 127516 66666
rect 127460 66612 127516 66614
rect 127564 66666 127620 66668
rect 127564 66614 127566 66666
rect 127566 66614 127618 66666
rect 127618 66614 127620 66666
rect 127564 66612 127620 66614
rect 127356 65098 127412 65100
rect 127356 65046 127358 65098
rect 127358 65046 127410 65098
rect 127410 65046 127412 65098
rect 127356 65044 127412 65046
rect 127460 65098 127516 65100
rect 127460 65046 127462 65098
rect 127462 65046 127514 65098
rect 127514 65046 127516 65098
rect 127460 65044 127516 65046
rect 127564 65098 127620 65100
rect 127564 65046 127566 65098
rect 127566 65046 127618 65098
rect 127618 65046 127620 65098
rect 127564 65044 127620 65046
rect 127356 63530 127412 63532
rect 127356 63478 127358 63530
rect 127358 63478 127410 63530
rect 127410 63478 127412 63530
rect 127356 63476 127412 63478
rect 127460 63530 127516 63532
rect 127460 63478 127462 63530
rect 127462 63478 127514 63530
rect 127514 63478 127516 63530
rect 127460 63476 127516 63478
rect 127564 63530 127620 63532
rect 127564 63478 127566 63530
rect 127566 63478 127618 63530
rect 127618 63478 127620 63530
rect 127564 63476 127620 63478
rect 127356 61962 127412 61964
rect 127356 61910 127358 61962
rect 127358 61910 127410 61962
rect 127410 61910 127412 61962
rect 127356 61908 127412 61910
rect 127460 61962 127516 61964
rect 127460 61910 127462 61962
rect 127462 61910 127514 61962
rect 127514 61910 127516 61962
rect 127460 61908 127516 61910
rect 127564 61962 127620 61964
rect 127564 61910 127566 61962
rect 127566 61910 127618 61962
rect 127618 61910 127620 61962
rect 127564 61908 127620 61910
rect 127356 60394 127412 60396
rect 127356 60342 127358 60394
rect 127358 60342 127410 60394
rect 127410 60342 127412 60394
rect 127356 60340 127412 60342
rect 127460 60394 127516 60396
rect 127460 60342 127462 60394
rect 127462 60342 127514 60394
rect 127514 60342 127516 60394
rect 127460 60340 127516 60342
rect 127564 60394 127620 60396
rect 127564 60342 127566 60394
rect 127566 60342 127618 60394
rect 127618 60342 127620 60394
rect 127564 60340 127620 60342
rect 127356 58826 127412 58828
rect 127356 58774 127358 58826
rect 127358 58774 127410 58826
rect 127410 58774 127412 58826
rect 127356 58772 127412 58774
rect 127460 58826 127516 58828
rect 127460 58774 127462 58826
rect 127462 58774 127514 58826
rect 127514 58774 127516 58826
rect 127460 58772 127516 58774
rect 127564 58826 127620 58828
rect 127564 58774 127566 58826
rect 127566 58774 127618 58826
rect 127618 58774 127620 58826
rect 127564 58772 127620 58774
rect 127356 57258 127412 57260
rect 127356 57206 127358 57258
rect 127358 57206 127410 57258
rect 127410 57206 127412 57258
rect 127356 57204 127412 57206
rect 127460 57258 127516 57260
rect 127460 57206 127462 57258
rect 127462 57206 127514 57258
rect 127514 57206 127516 57258
rect 127460 57204 127516 57206
rect 127564 57258 127620 57260
rect 127564 57206 127566 57258
rect 127566 57206 127618 57258
rect 127618 57206 127620 57258
rect 127564 57204 127620 57206
rect 127356 55690 127412 55692
rect 127356 55638 127358 55690
rect 127358 55638 127410 55690
rect 127410 55638 127412 55690
rect 127356 55636 127412 55638
rect 127460 55690 127516 55692
rect 127460 55638 127462 55690
rect 127462 55638 127514 55690
rect 127514 55638 127516 55690
rect 127460 55636 127516 55638
rect 127564 55690 127620 55692
rect 127564 55638 127566 55690
rect 127566 55638 127618 55690
rect 127618 55638 127620 55690
rect 127564 55636 127620 55638
rect 127356 54122 127412 54124
rect 127356 54070 127358 54122
rect 127358 54070 127410 54122
rect 127410 54070 127412 54122
rect 127356 54068 127412 54070
rect 127460 54122 127516 54124
rect 127460 54070 127462 54122
rect 127462 54070 127514 54122
rect 127514 54070 127516 54122
rect 127460 54068 127516 54070
rect 127564 54122 127620 54124
rect 127564 54070 127566 54122
rect 127566 54070 127618 54122
rect 127618 54070 127620 54122
rect 127564 54068 127620 54070
rect 127356 52554 127412 52556
rect 127356 52502 127358 52554
rect 127358 52502 127410 52554
rect 127410 52502 127412 52554
rect 127356 52500 127412 52502
rect 127460 52554 127516 52556
rect 127460 52502 127462 52554
rect 127462 52502 127514 52554
rect 127514 52502 127516 52554
rect 127460 52500 127516 52502
rect 127564 52554 127620 52556
rect 127564 52502 127566 52554
rect 127566 52502 127618 52554
rect 127618 52502 127620 52554
rect 127564 52500 127620 52502
rect 127356 50986 127412 50988
rect 127356 50934 127358 50986
rect 127358 50934 127410 50986
rect 127410 50934 127412 50986
rect 127356 50932 127412 50934
rect 127460 50986 127516 50988
rect 127460 50934 127462 50986
rect 127462 50934 127514 50986
rect 127514 50934 127516 50986
rect 127460 50932 127516 50934
rect 127564 50986 127620 50988
rect 127564 50934 127566 50986
rect 127566 50934 127618 50986
rect 127618 50934 127620 50986
rect 127564 50932 127620 50934
rect 127356 49418 127412 49420
rect 127356 49366 127358 49418
rect 127358 49366 127410 49418
rect 127410 49366 127412 49418
rect 127356 49364 127412 49366
rect 127460 49418 127516 49420
rect 127460 49366 127462 49418
rect 127462 49366 127514 49418
rect 127514 49366 127516 49418
rect 127460 49364 127516 49366
rect 127564 49418 127620 49420
rect 127564 49366 127566 49418
rect 127566 49366 127618 49418
rect 127618 49366 127620 49418
rect 127564 49364 127620 49366
rect 127356 47850 127412 47852
rect 127356 47798 127358 47850
rect 127358 47798 127410 47850
rect 127410 47798 127412 47850
rect 127356 47796 127412 47798
rect 127460 47850 127516 47852
rect 127460 47798 127462 47850
rect 127462 47798 127514 47850
rect 127514 47798 127516 47850
rect 127460 47796 127516 47798
rect 127564 47850 127620 47852
rect 127564 47798 127566 47850
rect 127566 47798 127618 47850
rect 127618 47798 127620 47850
rect 127564 47796 127620 47798
rect 127356 46282 127412 46284
rect 127356 46230 127358 46282
rect 127358 46230 127410 46282
rect 127410 46230 127412 46282
rect 127356 46228 127412 46230
rect 127460 46282 127516 46284
rect 127460 46230 127462 46282
rect 127462 46230 127514 46282
rect 127514 46230 127516 46282
rect 127460 46228 127516 46230
rect 127564 46282 127620 46284
rect 127564 46230 127566 46282
rect 127566 46230 127618 46282
rect 127618 46230 127620 46282
rect 127564 46228 127620 46230
rect 127356 44714 127412 44716
rect 127356 44662 127358 44714
rect 127358 44662 127410 44714
rect 127410 44662 127412 44714
rect 127356 44660 127412 44662
rect 127460 44714 127516 44716
rect 127460 44662 127462 44714
rect 127462 44662 127514 44714
rect 127514 44662 127516 44714
rect 127460 44660 127516 44662
rect 127564 44714 127620 44716
rect 127564 44662 127566 44714
rect 127566 44662 127618 44714
rect 127618 44662 127620 44714
rect 127564 44660 127620 44662
rect 127356 43146 127412 43148
rect 127356 43094 127358 43146
rect 127358 43094 127410 43146
rect 127410 43094 127412 43146
rect 127356 43092 127412 43094
rect 127460 43146 127516 43148
rect 127460 43094 127462 43146
rect 127462 43094 127514 43146
rect 127514 43094 127516 43146
rect 127460 43092 127516 43094
rect 127564 43146 127620 43148
rect 127564 43094 127566 43146
rect 127566 43094 127618 43146
rect 127618 43094 127620 43146
rect 127564 43092 127620 43094
rect 127356 41578 127412 41580
rect 127356 41526 127358 41578
rect 127358 41526 127410 41578
rect 127410 41526 127412 41578
rect 127356 41524 127412 41526
rect 127460 41578 127516 41580
rect 127460 41526 127462 41578
rect 127462 41526 127514 41578
rect 127514 41526 127516 41578
rect 127460 41524 127516 41526
rect 127564 41578 127620 41580
rect 127564 41526 127566 41578
rect 127566 41526 127618 41578
rect 127618 41526 127620 41578
rect 127564 41524 127620 41526
rect 127356 40010 127412 40012
rect 127356 39958 127358 40010
rect 127358 39958 127410 40010
rect 127410 39958 127412 40010
rect 127356 39956 127412 39958
rect 127460 40010 127516 40012
rect 127460 39958 127462 40010
rect 127462 39958 127514 40010
rect 127514 39958 127516 40010
rect 127460 39956 127516 39958
rect 127564 40010 127620 40012
rect 127564 39958 127566 40010
rect 127566 39958 127618 40010
rect 127618 39958 127620 40010
rect 127564 39956 127620 39958
rect 127356 38442 127412 38444
rect 127356 38390 127358 38442
rect 127358 38390 127410 38442
rect 127410 38390 127412 38442
rect 127356 38388 127412 38390
rect 127460 38442 127516 38444
rect 127460 38390 127462 38442
rect 127462 38390 127514 38442
rect 127514 38390 127516 38442
rect 127460 38388 127516 38390
rect 127564 38442 127620 38444
rect 127564 38390 127566 38442
rect 127566 38390 127618 38442
rect 127618 38390 127620 38442
rect 127564 38388 127620 38390
rect 127356 36874 127412 36876
rect 127356 36822 127358 36874
rect 127358 36822 127410 36874
rect 127410 36822 127412 36874
rect 127356 36820 127412 36822
rect 127460 36874 127516 36876
rect 127460 36822 127462 36874
rect 127462 36822 127514 36874
rect 127514 36822 127516 36874
rect 127460 36820 127516 36822
rect 127564 36874 127620 36876
rect 127564 36822 127566 36874
rect 127566 36822 127618 36874
rect 127618 36822 127620 36874
rect 127564 36820 127620 36822
rect 127356 35306 127412 35308
rect 127356 35254 127358 35306
rect 127358 35254 127410 35306
rect 127410 35254 127412 35306
rect 127356 35252 127412 35254
rect 127460 35306 127516 35308
rect 127460 35254 127462 35306
rect 127462 35254 127514 35306
rect 127514 35254 127516 35306
rect 127460 35252 127516 35254
rect 127564 35306 127620 35308
rect 127564 35254 127566 35306
rect 127566 35254 127618 35306
rect 127618 35254 127620 35306
rect 127564 35252 127620 35254
rect 127356 33738 127412 33740
rect 127356 33686 127358 33738
rect 127358 33686 127410 33738
rect 127410 33686 127412 33738
rect 127356 33684 127412 33686
rect 127460 33738 127516 33740
rect 127460 33686 127462 33738
rect 127462 33686 127514 33738
rect 127514 33686 127516 33738
rect 127460 33684 127516 33686
rect 127564 33738 127620 33740
rect 127564 33686 127566 33738
rect 127566 33686 127618 33738
rect 127618 33686 127620 33738
rect 127564 33684 127620 33686
rect 127356 32170 127412 32172
rect 127356 32118 127358 32170
rect 127358 32118 127410 32170
rect 127410 32118 127412 32170
rect 127356 32116 127412 32118
rect 127460 32170 127516 32172
rect 127460 32118 127462 32170
rect 127462 32118 127514 32170
rect 127514 32118 127516 32170
rect 127460 32116 127516 32118
rect 127564 32170 127620 32172
rect 127564 32118 127566 32170
rect 127566 32118 127618 32170
rect 127618 32118 127620 32170
rect 127564 32116 127620 32118
rect 127356 30602 127412 30604
rect 127356 30550 127358 30602
rect 127358 30550 127410 30602
rect 127410 30550 127412 30602
rect 127356 30548 127412 30550
rect 127460 30602 127516 30604
rect 127460 30550 127462 30602
rect 127462 30550 127514 30602
rect 127514 30550 127516 30602
rect 127460 30548 127516 30550
rect 127564 30602 127620 30604
rect 127564 30550 127566 30602
rect 127566 30550 127618 30602
rect 127618 30550 127620 30602
rect 127564 30548 127620 30550
rect 127356 29034 127412 29036
rect 127356 28982 127358 29034
rect 127358 28982 127410 29034
rect 127410 28982 127412 29034
rect 127356 28980 127412 28982
rect 127460 29034 127516 29036
rect 127460 28982 127462 29034
rect 127462 28982 127514 29034
rect 127514 28982 127516 29034
rect 127460 28980 127516 28982
rect 127564 29034 127620 29036
rect 127564 28982 127566 29034
rect 127566 28982 127618 29034
rect 127618 28982 127620 29034
rect 127564 28980 127620 28982
rect 126364 28588 126420 28644
rect 125244 9884 125300 9940
rect 125692 19180 125748 19236
rect 124796 6300 124852 6356
rect 124348 3500 124404 3556
rect 124236 3330 124292 3332
rect 124236 3278 124238 3330
rect 124238 3278 124290 3330
rect 124290 3278 124292 3330
rect 124236 3276 124292 3278
rect 125020 5740 125076 5796
rect 125020 5180 125076 5236
rect 124908 5122 124964 5124
rect 124908 5070 124910 5122
rect 124910 5070 124962 5122
rect 124962 5070 124964 5122
rect 124908 5068 124964 5070
rect 124796 4172 124852 4228
rect 125132 4956 125188 5012
rect 125692 6636 125748 6692
rect 125916 6636 125972 6692
rect 125356 5964 125412 6020
rect 125356 5122 125412 5124
rect 125356 5070 125358 5122
rect 125358 5070 125410 5122
rect 125410 5070 125412 5122
rect 125356 5068 125412 5070
rect 125132 4060 125188 4116
rect 125580 5794 125636 5796
rect 125580 5742 125582 5794
rect 125582 5742 125634 5794
rect 125634 5742 125636 5794
rect 125580 5740 125636 5742
rect 125580 5404 125636 5460
rect 125356 3612 125412 3668
rect 125244 3500 125300 3556
rect 125132 3164 125188 3220
rect 124908 2940 124964 2996
rect 125804 5964 125860 6020
rect 125804 5516 125860 5572
rect 125916 5404 125972 5460
rect 126028 5234 126084 5236
rect 126028 5182 126030 5234
rect 126030 5182 126082 5234
rect 126082 5182 126084 5234
rect 126028 5180 126084 5182
rect 125804 4450 125860 4452
rect 125804 4398 125806 4450
rect 125806 4398 125858 4450
rect 125858 4398 125860 4450
rect 125804 4396 125860 4398
rect 125692 4172 125748 4228
rect 125580 3276 125636 3332
rect 125804 3612 125860 3668
rect 126140 3836 126196 3892
rect 127356 27466 127412 27468
rect 127356 27414 127358 27466
rect 127358 27414 127410 27466
rect 127410 27414 127412 27466
rect 127356 27412 127412 27414
rect 127460 27466 127516 27468
rect 127460 27414 127462 27466
rect 127462 27414 127514 27466
rect 127514 27414 127516 27466
rect 127460 27412 127516 27414
rect 127564 27466 127620 27468
rect 127564 27414 127566 27466
rect 127566 27414 127618 27466
rect 127618 27414 127620 27466
rect 127564 27412 127620 27414
rect 127356 25898 127412 25900
rect 127356 25846 127358 25898
rect 127358 25846 127410 25898
rect 127410 25846 127412 25898
rect 127356 25844 127412 25846
rect 127460 25898 127516 25900
rect 127460 25846 127462 25898
rect 127462 25846 127514 25898
rect 127514 25846 127516 25898
rect 127460 25844 127516 25846
rect 127564 25898 127620 25900
rect 127564 25846 127566 25898
rect 127566 25846 127618 25898
rect 127618 25846 127620 25898
rect 127564 25844 127620 25846
rect 127356 24330 127412 24332
rect 127356 24278 127358 24330
rect 127358 24278 127410 24330
rect 127410 24278 127412 24330
rect 127356 24276 127412 24278
rect 127460 24330 127516 24332
rect 127460 24278 127462 24330
rect 127462 24278 127514 24330
rect 127514 24278 127516 24330
rect 127460 24276 127516 24278
rect 127564 24330 127620 24332
rect 127564 24278 127566 24330
rect 127566 24278 127618 24330
rect 127618 24278 127620 24330
rect 127564 24276 127620 24278
rect 127356 22762 127412 22764
rect 127356 22710 127358 22762
rect 127358 22710 127410 22762
rect 127410 22710 127412 22762
rect 127356 22708 127412 22710
rect 127460 22762 127516 22764
rect 127460 22710 127462 22762
rect 127462 22710 127514 22762
rect 127514 22710 127516 22762
rect 127460 22708 127516 22710
rect 127564 22762 127620 22764
rect 127564 22710 127566 22762
rect 127566 22710 127618 22762
rect 127618 22710 127620 22762
rect 127564 22708 127620 22710
rect 130396 22092 130452 22148
rect 127356 21194 127412 21196
rect 127356 21142 127358 21194
rect 127358 21142 127410 21194
rect 127410 21142 127412 21194
rect 127356 21140 127412 21142
rect 127460 21194 127516 21196
rect 127460 21142 127462 21194
rect 127462 21142 127514 21194
rect 127514 21142 127516 21194
rect 127460 21140 127516 21142
rect 127564 21194 127620 21196
rect 127564 21142 127566 21194
rect 127566 21142 127618 21194
rect 127618 21142 127620 21194
rect 127564 21140 127620 21142
rect 127148 20636 127204 20692
rect 126476 5964 126532 6020
rect 126924 6690 126980 6692
rect 126924 6638 126926 6690
rect 126926 6638 126978 6690
rect 126978 6638 126980 6690
rect 126924 6636 126980 6638
rect 128492 20188 128548 20244
rect 127356 19626 127412 19628
rect 127356 19574 127358 19626
rect 127358 19574 127410 19626
rect 127410 19574 127412 19626
rect 127356 19572 127412 19574
rect 127460 19626 127516 19628
rect 127460 19574 127462 19626
rect 127462 19574 127514 19626
rect 127514 19574 127516 19626
rect 127460 19572 127516 19574
rect 127564 19626 127620 19628
rect 127564 19574 127566 19626
rect 127566 19574 127618 19626
rect 127618 19574 127620 19626
rect 127564 19572 127620 19574
rect 127356 18058 127412 18060
rect 127356 18006 127358 18058
rect 127358 18006 127410 18058
rect 127410 18006 127412 18058
rect 127356 18004 127412 18006
rect 127460 18058 127516 18060
rect 127460 18006 127462 18058
rect 127462 18006 127514 18058
rect 127514 18006 127516 18058
rect 127460 18004 127516 18006
rect 127564 18058 127620 18060
rect 127564 18006 127566 18058
rect 127566 18006 127618 18058
rect 127618 18006 127620 18058
rect 127564 18004 127620 18006
rect 127356 16490 127412 16492
rect 127356 16438 127358 16490
rect 127358 16438 127410 16490
rect 127410 16438 127412 16490
rect 127356 16436 127412 16438
rect 127460 16490 127516 16492
rect 127460 16438 127462 16490
rect 127462 16438 127514 16490
rect 127514 16438 127516 16490
rect 127460 16436 127516 16438
rect 127564 16490 127620 16492
rect 127564 16438 127566 16490
rect 127566 16438 127618 16490
rect 127618 16438 127620 16490
rect 127564 16436 127620 16438
rect 127356 14922 127412 14924
rect 127356 14870 127358 14922
rect 127358 14870 127410 14922
rect 127410 14870 127412 14922
rect 127356 14868 127412 14870
rect 127460 14922 127516 14924
rect 127460 14870 127462 14922
rect 127462 14870 127514 14922
rect 127514 14870 127516 14922
rect 127460 14868 127516 14870
rect 127564 14922 127620 14924
rect 127564 14870 127566 14922
rect 127566 14870 127618 14922
rect 127618 14870 127620 14922
rect 127564 14868 127620 14870
rect 127356 13354 127412 13356
rect 127356 13302 127358 13354
rect 127358 13302 127410 13354
rect 127410 13302 127412 13354
rect 127356 13300 127412 13302
rect 127460 13354 127516 13356
rect 127460 13302 127462 13354
rect 127462 13302 127514 13354
rect 127514 13302 127516 13354
rect 127460 13300 127516 13302
rect 127564 13354 127620 13356
rect 127564 13302 127566 13354
rect 127566 13302 127618 13354
rect 127618 13302 127620 13354
rect 127564 13300 127620 13302
rect 127356 11786 127412 11788
rect 127356 11734 127358 11786
rect 127358 11734 127410 11786
rect 127410 11734 127412 11786
rect 127356 11732 127412 11734
rect 127460 11786 127516 11788
rect 127460 11734 127462 11786
rect 127462 11734 127514 11786
rect 127514 11734 127516 11786
rect 127460 11732 127516 11734
rect 127564 11786 127620 11788
rect 127564 11734 127566 11786
rect 127566 11734 127618 11786
rect 127618 11734 127620 11786
rect 127564 11732 127620 11734
rect 128044 11452 128100 11508
rect 127356 10218 127412 10220
rect 127356 10166 127358 10218
rect 127358 10166 127410 10218
rect 127410 10166 127412 10218
rect 127356 10164 127412 10166
rect 127460 10218 127516 10220
rect 127460 10166 127462 10218
rect 127462 10166 127514 10218
rect 127514 10166 127516 10218
rect 127460 10164 127516 10166
rect 127564 10218 127620 10220
rect 127564 10166 127566 10218
rect 127566 10166 127618 10218
rect 127618 10166 127620 10218
rect 127564 10164 127620 10166
rect 127356 8650 127412 8652
rect 127356 8598 127358 8650
rect 127358 8598 127410 8650
rect 127410 8598 127412 8650
rect 127356 8596 127412 8598
rect 127460 8650 127516 8652
rect 127460 8598 127462 8650
rect 127462 8598 127514 8650
rect 127514 8598 127516 8650
rect 127460 8596 127516 8598
rect 127564 8650 127620 8652
rect 127564 8598 127566 8650
rect 127566 8598 127618 8650
rect 127618 8598 127620 8650
rect 127564 8596 127620 8598
rect 127356 7082 127412 7084
rect 127356 7030 127358 7082
rect 127358 7030 127410 7082
rect 127410 7030 127412 7082
rect 127356 7028 127412 7030
rect 127460 7082 127516 7084
rect 127460 7030 127462 7082
rect 127462 7030 127514 7082
rect 127514 7030 127516 7082
rect 127460 7028 127516 7030
rect 127564 7082 127620 7084
rect 127564 7030 127566 7082
rect 127566 7030 127618 7082
rect 127618 7030 127620 7082
rect 127564 7028 127620 7030
rect 127820 6524 127876 6580
rect 126812 5794 126868 5796
rect 126812 5742 126814 5794
rect 126814 5742 126866 5794
rect 126866 5742 126868 5794
rect 126812 5740 126868 5742
rect 126252 4284 126308 4340
rect 126028 3330 126084 3332
rect 126028 3278 126030 3330
rect 126030 3278 126082 3330
rect 126082 3278 126084 3330
rect 126028 3276 126084 3278
rect 126140 2828 126196 2884
rect 126364 3388 126420 3444
rect 126812 4508 126868 4564
rect 126700 3836 126756 3892
rect 126252 1148 126308 1204
rect 127708 5852 127764 5908
rect 127356 5514 127412 5516
rect 127356 5462 127358 5514
rect 127358 5462 127410 5514
rect 127410 5462 127412 5514
rect 127356 5460 127412 5462
rect 127460 5514 127516 5516
rect 127460 5462 127462 5514
rect 127462 5462 127514 5514
rect 127514 5462 127516 5514
rect 127460 5460 127516 5462
rect 127564 5514 127620 5516
rect 127564 5462 127566 5514
rect 127566 5462 127618 5514
rect 127618 5462 127620 5514
rect 127708 5516 127764 5572
rect 129836 12684 129892 12740
rect 129276 12012 129332 12068
rect 128492 10108 128548 10164
rect 129052 10108 129108 10164
rect 128604 7532 128660 7588
rect 128044 6412 128100 6468
rect 128156 6748 128212 6804
rect 127932 5964 127988 6020
rect 128268 5906 128324 5908
rect 128268 5854 128270 5906
rect 128270 5854 128322 5906
rect 128322 5854 128324 5906
rect 128268 5852 128324 5854
rect 127564 5460 127620 5462
rect 128604 6748 128660 6804
rect 127148 5180 127204 5236
rect 128492 6412 128548 6468
rect 127260 5122 127316 5124
rect 127260 5070 127262 5122
rect 127262 5070 127314 5122
rect 127314 5070 127316 5122
rect 127260 5068 127316 5070
rect 127596 5068 127652 5124
rect 127708 4956 127764 5012
rect 127036 3500 127092 3556
rect 126812 1484 126868 1540
rect 126924 3388 126980 3444
rect 127356 3946 127412 3948
rect 127356 3894 127358 3946
rect 127358 3894 127410 3946
rect 127410 3894 127412 3946
rect 127356 3892 127412 3894
rect 127460 3946 127516 3948
rect 127460 3894 127462 3946
rect 127462 3894 127514 3946
rect 127514 3894 127516 3946
rect 127460 3892 127516 3894
rect 127564 3946 127620 3948
rect 127564 3894 127566 3946
rect 127566 3894 127618 3946
rect 127618 3894 127620 3946
rect 127564 3892 127620 3894
rect 127596 3724 127652 3780
rect 127260 3554 127316 3556
rect 127260 3502 127262 3554
rect 127262 3502 127314 3554
rect 127314 3502 127316 3554
rect 127260 3500 127316 3502
rect 127484 3500 127540 3556
rect 127036 3052 127092 3108
rect 127932 4562 127988 4564
rect 127932 4510 127934 4562
rect 127934 4510 127986 4562
rect 127986 4510 127988 4562
rect 127932 4508 127988 4510
rect 128156 5122 128212 5124
rect 128156 5070 128158 5122
rect 128158 5070 128210 5122
rect 128210 5070 128212 5122
rect 128156 5068 128212 5070
rect 128492 5068 128548 5124
rect 128604 5964 128660 6020
rect 128044 4284 128100 4340
rect 128156 4844 128212 4900
rect 128716 4284 128772 4340
rect 128940 6860 128996 6916
rect 129276 7644 129332 7700
rect 129052 4450 129108 4452
rect 129052 4398 129054 4450
rect 129054 4398 129106 4450
rect 129106 4398 129108 4450
rect 129052 4396 129108 4398
rect 129276 5906 129332 5908
rect 129276 5854 129278 5906
rect 129278 5854 129330 5906
rect 129330 5854 129332 5906
rect 129276 5852 129332 5854
rect 129276 4620 129332 4676
rect 128044 3836 128100 3892
rect 127820 3164 127876 3220
rect 127820 2268 127876 2324
rect 128492 3612 128548 3668
rect 128604 3948 128660 4004
rect 128156 3330 128212 3332
rect 128156 3278 128158 3330
rect 128158 3278 128210 3330
rect 128210 3278 128212 3330
rect 128156 3276 128212 3278
rect 129164 4060 129220 4116
rect 129164 3612 129220 3668
rect 128940 3388 128996 3444
rect 129612 5964 129668 6020
rect 130172 7980 130228 8036
rect 129948 7698 130004 7700
rect 129948 7646 129950 7698
rect 129950 7646 130002 7698
rect 130002 7646 130004 7698
rect 129948 7644 130004 7646
rect 130060 7420 130116 7476
rect 130060 6412 130116 6468
rect 129724 4620 129780 4676
rect 129948 4844 130004 4900
rect 130060 5404 130116 5460
rect 129836 3836 129892 3892
rect 130284 7644 130340 7700
rect 130396 7474 130452 7476
rect 130396 7422 130398 7474
rect 130398 7422 130450 7474
rect 130450 7422 130452 7474
rect 130396 7420 130452 7422
rect 144060 117180 144116 117236
rect 144956 117180 145012 117236
rect 148764 116620 148820 116676
rect 149548 116620 149604 116676
rect 145628 116508 145684 116564
rect 147532 116562 147588 116564
rect 147532 116510 147534 116562
rect 147534 116510 147586 116562
rect 147586 116510 147588 116562
rect 147532 116508 147588 116510
rect 153468 116956 153524 117012
rect 150332 116508 150388 116564
rect 151452 116562 151508 116564
rect 151452 116510 151454 116562
rect 151454 116510 151506 116562
rect 151506 116510 151508 116562
rect 151452 116508 151508 116510
rect 142716 116058 142772 116060
rect 142716 116006 142718 116058
rect 142718 116006 142770 116058
rect 142770 116006 142772 116058
rect 142716 116004 142772 116006
rect 142820 116058 142876 116060
rect 142820 116006 142822 116058
rect 142822 116006 142874 116058
rect 142874 116006 142876 116058
rect 142820 116004 142876 116006
rect 142924 116058 142980 116060
rect 142924 116006 142926 116058
rect 142926 116006 142978 116058
rect 142978 116006 142980 116058
rect 142924 116004 142980 116006
rect 146076 116450 146132 116452
rect 146076 116398 146078 116450
rect 146078 116398 146130 116450
rect 146130 116398 146132 116450
rect 146076 116396 146132 116398
rect 146860 116450 146916 116452
rect 146860 116398 146862 116450
rect 146862 116398 146914 116450
rect 146914 116398 146916 116450
rect 146860 116396 146916 116398
rect 153468 116396 153524 116452
rect 140924 115724 140980 115780
rect 142044 115778 142100 115780
rect 142044 115726 142046 115778
rect 142046 115726 142098 115778
rect 142098 115726 142100 115778
rect 142044 115724 142100 115726
rect 138460 115666 138516 115668
rect 138460 115614 138462 115666
rect 138462 115614 138514 115666
rect 138514 115614 138516 115666
rect 138460 115612 138516 115614
rect 139132 115666 139188 115668
rect 139132 115614 139134 115666
rect 139134 115614 139186 115666
rect 139186 115614 139188 115666
rect 139132 115612 139188 115614
rect 133980 23884 134036 23940
rect 131740 16716 131796 16772
rect 133532 22316 133588 22372
rect 131516 15484 131572 15540
rect 130732 10556 130788 10612
rect 130620 8034 130676 8036
rect 130620 7982 130622 8034
rect 130622 7982 130674 8034
rect 130674 7982 130676 8034
rect 130620 7980 130676 7982
rect 130620 6690 130676 6692
rect 130620 6638 130622 6690
rect 130622 6638 130674 6690
rect 130674 6638 130676 6690
rect 130620 6636 130676 6638
rect 130508 6524 130564 6580
rect 131068 8034 131124 8036
rect 131068 7982 131070 8034
rect 131070 7982 131122 8034
rect 131122 7982 131124 8034
rect 131068 7980 131124 7982
rect 130844 7698 130900 7700
rect 130844 7646 130846 7698
rect 130846 7646 130898 7698
rect 130898 7646 130900 7698
rect 130844 7644 130900 7646
rect 130956 6860 131012 6916
rect 130844 6636 130900 6692
rect 130060 3724 130116 3780
rect 130284 3836 130340 3892
rect 130172 3442 130228 3444
rect 130172 3390 130174 3442
rect 130174 3390 130226 3442
rect 130226 3390 130228 3442
rect 130172 3388 130228 3390
rect 129500 3164 129556 3220
rect 129388 1036 129444 1092
rect 130060 3164 130116 3220
rect 130620 5010 130676 5012
rect 130620 4958 130622 5010
rect 130622 4958 130674 5010
rect 130674 4958 130676 5010
rect 130620 4956 130676 4958
rect 130508 2716 130564 2772
rect 130844 4844 130900 4900
rect 130844 4620 130900 4676
rect 130732 2268 130788 2324
rect 130844 3500 130900 3556
rect 98588 700 98644 756
rect 131180 6076 131236 6132
rect 131180 5068 131236 5124
rect 131068 4732 131124 4788
rect 131068 4450 131124 4452
rect 131068 4398 131070 4450
rect 131070 4398 131122 4450
rect 131122 4398 131124 4450
rect 131068 4396 131124 4398
rect 131964 7474 132020 7476
rect 131964 7422 131966 7474
rect 131966 7422 132018 7474
rect 132018 7422 132020 7474
rect 131964 7420 132020 7422
rect 131740 6018 131796 6020
rect 131740 5966 131742 6018
rect 131742 5966 131794 6018
rect 131794 5966 131796 6018
rect 131740 5964 131796 5966
rect 132076 5628 132132 5684
rect 131292 3612 131348 3668
rect 131740 5234 131796 5236
rect 131740 5182 131742 5234
rect 131742 5182 131794 5234
rect 131794 5182 131796 5234
rect 131740 5180 131796 5182
rect 130956 3388 131012 3444
rect 131180 2492 131236 2548
rect 131628 4508 131684 4564
rect 131516 3612 131572 3668
rect 131852 3276 131908 3332
rect 132412 7698 132468 7700
rect 132412 7646 132414 7698
rect 132414 7646 132466 7698
rect 132466 7646 132468 7698
rect 132412 7644 132468 7646
rect 132300 6860 132356 6916
rect 132636 6300 132692 6356
rect 132748 5292 132804 5348
rect 132188 3948 132244 4004
rect 132412 4284 132468 4340
rect 132188 3612 132244 3668
rect 131964 3164 132020 3220
rect 132972 6188 133028 6244
rect 133084 7644 133140 7700
rect 132972 6018 133028 6020
rect 132972 5966 132974 6018
rect 132974 5966 133026 6018
rect 133026 5966 133028 6018
rect 132972 5964 133028 5966
rect 133756 13468 133812 13524
rect 133532 7644 133588 7700
rect 133196 6188 133252 6244
rect 133196 5628 133252 5684
rect 133084 4620 133140 4676
rect 132636 3836 132692 3892
rect 133420 5346 133476 5348
rect 133420 5294 133422 5346
rect 133422 5294 133474 5346
rect 133474 5294 133476 5346
rect 133420 5292 133476 5294
rect 133868 6466 133924 6468
rect 133868 6414 133870 6466
rect 133870 6414 133922 6466
rect 133922 6414 133924 6466
rect 133868 6412 133924 6414
rect 135548 22428 135604 22484
rect 134764 18620 134820 18676
rect 134428 7698 134484 7700
rect 134428 7646 134430 7698
rect 134430 7646 134482 7698
rect 134482 7646 134484 7698
rect 134428 7644 134484 7646
rect 133980 5682 134036 5684
rect 133980 5630 133982 5682
rect 133982 5630 134034 5682
rect 134034 5630 134036 5682
rect 133980 5628 134036 5630
rect 133868 5404 133924 5460
rect 133644 5122 133700 5124
rect 133644 5070 133646 5122
rect 133646 5070 133698 5122
rect 133698 5070 133700 5122
rect 133644 5068 133700 5070
rect 133868 4956 133924 5012
rect 134652 7084 134708 7140
rect 133980 5068 134036 5124
rect 134204 6300 134260 6356
rect 133420 3724 133476 3780
rect 132524 3388 132580 3444
rect 132972 2604 133028 2660
rect 133756 4844 133812 4900
rect 133868 4732 133924 4788
rect 133756 4620 133812 4676
rect 134764 6636 134820 6692
rect 135548 7756 135604 7812
rect 134540 6018 134596 6020
rect 134540 5966 134542 6018
rect 134542 5966 134594 6018
rect 134594 5966 134596 6018
rect 134540 5964 134596 5966
rect 134540 5628 134596 5684
rect 134876 5906 134932 5908
rect 134876 5854 134878 5906
rect 134878 5854 134930 5906
rect 134930 5854 134932 5906
rect 134876 5852 134932 5854
rect 134764 5516 134820 5572
rect 134540 5404 134596 5460
rect 133868 4172 133924 4228
rect 133644 3500 133700 3556
rect 133756 3724 133812 3780
rect 134428 4338 134484 4340
rect 134428 4286 134430 4338
rect 134430 4286 134482 4338
rect 134482 4286 134484 4338
rect 134428 4284 134484 4286
rect 134652 4732 134708 4788
rect 134316 3948 134372 4004
rect 134204 3554 134260 3556
rect 134204 3502 134206 3554
rect 134206 3502 134258 3554
rect 134258 3502 134260 3554
rect 134204 3500 134260 3502
rect 135100 4956 135156 5012
rect 135324 6076 135380 6132
rect 135772 19068 135828 19124
rect 136780 17724 136836 17780
rect 136668 12236 136724 12292
rect 143164 115666 143220 115668
rect 143164 115614 143166 115666
rect 143166 115614 143218 115666
rect 143218 115614 143220 115666
rect 143164 115612 143220 115614
rect 143836 115666 143892 115668
rect 143836 115614 143838 115666
rect 143838 115614 143890 115666
rect 143890 115614 143892 115666
rect 143836 115612 143892 115614
rect 147868 115666 147924 115668
rect 147868 115614 147870 115666
rect 147870 115614 147922 115666
rect 147922 115614 147924 115666
rect 147868 115612 147924 115614
rect 148540 115666 148596 115668
rect 148540 115614 148542 115666
rect 148542 115614 148594 115666
rect 148594 115614 148596 115666
rect 148540 115612 148596 115614
rect 142716 114490 142772 114492
rect 142716 114438 142718 114490
rect 142718 114438 142770 114490
rect 142770 114438 142772 114490
rect 142716 114436 142772 114438
rect 142820 114490 142876 114492
rect 142820 114438 142822 114490
rect 142822 114438 142874 114490
rect 142874 114438 142876 114490
rect 142820 114436 142876 114438
rect 142924 114490 142980 114492
rect 142924 114438 142926 114490
rect 142926 114438 142978 114490
rect 142978 114438 142980 114490
rect 142924 114436 142980 114438
rect 142716 112922 142772 112924
rect 142716 112870 142718 112922
rect 142718 112870 142770 112922
rect 142770 112870 142772 112922
rect 142716 112868 142772 112870
rect 142820 112922 142876 112924
rect 142820 112870 142822 112922
rect 142822 112870 142874 112922
rect 142874 112870 142876 112922
rect 142820 112868 142876 112870
rect 142924 112922 142980 112924
rect 142924 112870 142926 112922
rect 142926 112870 142978 112922
rect 142978 112870 142980 112922
rect 142924 112868 142980 112870
rect 142716 111354 142772 111356
rect 142716 111302 142718 111354
rect 142718 111302 142770 111354
rect 142770 111302 142772 111354
rect 142716 111300 142772 111302
rect 142820 111354 142876 111356
rect 142820 111302 142822 111354
rect 142822 111302 142874 111354
rect 142874 111302 142876 111354
rect 142820 111300 142876 111302
rect 142924 111354 142980 111356
rect 142924 111302 142926 111354
rect 142926 111302 142978 111354
rect 142978 111302 142980 111354
rect 142924 111300 142980 111302
rect 142716 109786 142772 109788
rect 142716 109734 142718 109786
rect 142718 109734 142770 109786
rect 142770 109734 142772 109786
rect 142716 109732 142772 109734
rect 142820 109786 142876 109788
rect 142820 109734 142822 109786
rect 142822 109734 142874 109786
rect 142874 109734 142876 109786
rect 142820 109732 142876 109734
rect 142924 109786 142980 109788
rect 142924 109734 142926 109786
rect 142926 109734 142978 109786
rect 142978 109734 142980 109786
rect 142924 109732 142980 109734
rect 142716 108218 142772 108220
rect 142716 108166 142718 108218
rect 142718 108166 142770 108218
rect 142770 108166 142772 108218
rect 142716 108164 142772 108166
rect 142820 108218 142876 108220
rect 142820 108166 142822 108218
rect 142822 108166 142874 108218
rect 142874 108166 142876 108218
rect 142820 108164 142876 108166
rect 142924 108218 142980 108220
rect 142924 108166 142926 108218
rect 142926 108166 142978 108218
rect 142978 108166 142980 108218
rect 142924 108164 142980 108166
rect 142716 106650 142772 106652
rect 142716 106598 142718 106650
rect 142718 106598 142770 106650
rect 142770 106598 142772 106650
rect 142716 106596 142772 106598
rect 142820 106650 142876 106652
rect 142820 106598 142822 106650
rect 142822 106598 142874 106650
rect 142874 106598 142876 106650
rect 142820 106596 142876 106598
rect 142924 106650 142980 106652
rect 142924 106598 142926 106650
rect 142926 106598 142978 106650
rect 142978 106598 142980 106650
rect 142924 106596 142980 106598
rect 142716 105082 142772 105084
rect 142716 105030 142718 105082
rect 142718 105030 142770 105082
rect 142770 105030 142772 105082
rect 142716 105028 142772 105030
rect 142820 105082 142876 105084
rect 142820 105030 142822 105082
rect 142822 105030 142874 105082
rect 142874 105030 142876 105082
rect 142820 105028 142876 105030
rect 142924 105082 142980 105084
rect 142924 105030 142926 105082
rect 142926 105030 142978 105082
rect 142978 105030 142980 105082
rect 142924 105028 142980 105030
rect 142716 103514 142772 103516
rect 142716 103462 142718 103514
rect 142718 103462 142770 103514
rect 142770 103462 142772 103514
rect 142716 103460 142772 103462
rect 142820 103514 142876 103516
rect 142820 103462 142822 103514
rect 142822 103462 142874 103514
rect 142874 103462 142876 103514
rect 142820 103460 142876 103462
rect 142924 103514 142980 103516
rect 142924 103462 142926 103514
rect 142926 103462 142978 103514
rect 142978 103462 142980 103514
rect 142924 103460 142980 103462
rect 142716 101946 142772 101948
rect 142716 101894 142718 101946
rect 142718 101894 142770 101946
rect 142770 101894 142772 101946
rect 142716 101892 142772 101894
rect 142820 101946 142876 101948
rect 142820 101894 142822 101946
rect 142822 101894 142874 101946
rect 142874 101894 142876 101946
rect 142820 101892 142876 101894
rect 142924 101946 142980 101948
rect 142924 101894 142926 101946
rect 142926 101894 142978 101946
rect 142978 101894 142980 101946
rect 142924 101892 142980 101894
rect 142716 100378 142772 100380
rect 142716 100326 142718 100378
rect 142718 100326 142770 100378
rect 142770 100326 142772 100378
rect 142716 100324 142772 100326
rect 142820 100378 142876 100380
rect 142820 100326 142822 100378
rect 142822 100326 142874 100378
rect 142874 100326 142876 100378
rect 142820 100324 142876 100326
rect 142924 100378 142980 100380
rect 142924 100326 142926 100378
rect 142926 100326 142978 100378
rect 142978 100326 142980 100378
rect 142924 100324 142980 100326
rect 142716 98810 142772 98812
rect 142716 98758 142718 98810
rect 142718 98758 142770 98810
rect 142770 98758 142772 98810
rect 142716 98756 142772 98758
rect 142820 98810 142876 98812
rect 142820 98758 142822 98810
rect 142822 98758 142874 98810
rect 142874 98758 142876 98810
rect 142820 98756 142876 98758
rect 142924 98810 142980 98812
rect 142924 98758 142926 98810
rect 142926 98758 142978 98810
rect 142978 98758 142980 98810
rect 142924 98756 142980 98758
rect 142716 97242 142772 97244
rect 142716 97190 142718 97242
rect 142718 97190 142770 97242
rect 142770 97190 142772 97242
rect 142716 97188 142772 97190
rect 142820 97242 142876 97244
rect 142820 97190 142822 97242
rect 142822 97190 142874 97242
rect 142874 97190 142876 97242
rect 142820 97188 142876 97190
rect 142924 97242 142980 97244
rect 142924 97190 142926 97242
rect 142926 97190 142978 97242
rect 142978 97190 142980 97242
rect 142924 97188 142980 97190
rect 142716 95674 142772 95676
rect 142716 95622 142718 95674
rect 142718 95622 142770 95674
rect 142770 95622 142772 95674
rect 142716 95620 142772 95622
rect 142820 95674 142876 95676
rect 142820 95622 142822 95674
rect 142822 95622 142874 95674
rect 142874 95622 142876 95674
rect 142820 95620 142876 95622
rect 142924 95674 142980 95676
rect 142924 95622 142926 95674
rect 142926 95622 142978 95674
rect 142978 95622 142980 95674
rect 142924 95620 142980 95622
rect 142716 94106 142772 94108
rect 142716 94054 142718 94106
rect 142718 94054 142770 94106
rect 142770 94054 142772 94106
rect 142716 94052 142772 94054
rect 142820 94106 142876 94108
rect 142820 94054 142822 94106
rect 142822 94054 142874 94106
rect 142874 94054 142876 94106
rect 142820 94052 142876 94054
rect 142924 94106 142980 94108
rect 142924 94054 142926 94106
rect 142926 94054 142978 94106
rect 142978 94054 142980 94106
rect 142924 94052 142980 94054
rect 142716 92538 142772 92540
rect 142716 92486 142718 92538
rect 142718 92486 142770 92538
rect 142770 92486 142772 92538
rect 142716 92484 142772 92486
rect 142820 92538 142876 92540
rect 142820 92486 142822 92538
rect 142822 92486 142874 92538
rect 142874 92486 142876 92538
rect 142820 92484 142876 92486
rect 142924 92538 142980 92540
rect 142924 92486 142926 92538
rect 142926 92486 142978 92538
rect 142978 92486 142980 92538
rect 142924 92484 142980 92486
rect 142716 90970 142772 90972
rect 142716 90918 142718 90970
rect 142718 90918 142770 90970
rect 142770 90918 142772 90970
rect 142716 90916 142772 90918
rect 142820 90970 142876 90972
rect 142820 90918 142822 90970
rect 142822 90918 142874 90970
rect 142874 90918 142876 90970
rect 142820 90916 142876 90918
rect 142924 90970 142980 90972
rect 142924 90918 142926 90970
rect 142926 90918 142978 90970
rect 142978 90918 142980 90970
rect 142924 90916 142980 90918
rect 142716 89402 142772 89404
rect 142716 89350 142718 89402
rect 142718 89350 142770 89402
rect 142770 89350 142772 89402
rect 142716 89348 142772 89350
rect 142820 89402 142876 89404
rect 142820 89350 142822 89402
rect 142822 89350 142874 89402
rect 142874 89350 142876 89402
rect 142820 89348 142876 89350
rect 142924 89402 142980 89404
rect 142924 89350 142926 89402
rect 142926 89350 142978 89402
rect 142978 89350 142980 89402
rect 142924 89348 142980 89350
rect 142716 87834 142772 87836
rect 142716 87782 142718 87834
rect 142718 87782 142770 87834
rect 142770 87782 142772 87834
rect 142716 87780 142772 87782
rect 142820 87834 142876 87836
rect 142820 87782 142822 87834
rect 142822 87782 142874 87834
rect 142874 87782 142876 87834
rect 142820 87780 142876 87782
rect 142924 87834 142980 87836
rect 142924 87782 142926 87834
rect 142926 87782 142978 87834
rect 142978 87782 142980 87834
rect 142924 87780 142980 87782
rect 142716 86266 142772 86268
rect 142716 86214 142718 86266
rect 142718 86214 142770 86266
rect 142770 86214 142772 86266
rect 142716 86212 142772 86214
rect 142820 86266 142876 86268
rect 142820 86214 142822 86266
rect 142822 86214 142874 86266
rect 142874 86214 142876 86266
rect 142820 86212 142876 86214
rect 142924 86266 142980 86268
rect 142924 86214 142926 86266
rect 142926 86214 142978 86266
rect 142978 86214 142980 86266
rect 142924 86212 142980 86214
rect 142716 84698 142772 84700
rect 142716 84646 142718 84698
rect 142718 84646 142770 84698
rect 142770 84646 142772 84698
rect 142716 84644 142772 84646
rect 142820 84698 142876 84700
rect 142820 84646 142822 84698
rect 142822 84646 142874 84698
rect 142874 84646 142876 84698
rect 142820 84644 142876 84646
rect 142924 84698 142980 84700
rect 142924 84646 142926 84698
rect 142926 84646 142978 84698
rect 142978 84646 142980 84698
rect 142924 84644 142980 84646
rect 142716 83130 142772 83132
rect 142716 83078 142718 83130
rect 142718 83078 142770 83130
rect 142770 83078 142772 83130
rect 142716 83076 142772 83078
rect 142820 83130 142876 83132
rect 142820 83078 142822 83130
rect 142822 83078 142874 83130
rect 142874 83078 142876 83130
rect 142820 83076 142876 83078
rect 142924 83130 142980 83132
rect 142924 83078 142926 83130
rect 142926 83078 142978 83130
rect 142978 83078 142980 83130
rect 142924 83076 142980 83078
rect 142716 81562 142772 81564
rect 142716 81510 142718 81562
rect 142718 81510 142770 81562
rect 142770 81510 142772 81562
rect 142716 81508 142772 81510
rect 142820 81562 142876 81564
rect 142820 81510 142822 81562
rect 142822 81510 142874 81562
rect 142874 81510 142876 81562
rect 142820 81508 142876 81510
rect 142924 81562 142980 81564
rect 142924 81510 142926 81562
rect 142926 81510 142978 81562
rect 142978 81510 142980 81562
rect 142924 81508 142980 81510
rect 142716 79994 142772 79996
rect 142716 79942 142718 79994
rect 142718 79942 142770 79994
rect 142770 79942 142772 79994
rect 142716 79940 142772 79942
rect 142820 79994 142876 79996
rect 142820 79942 142822 79994
rect 142822 79942 142874 79994
rect 142874 79942 142876 79994
rect 142820 79940 142876 79942
rect 142924 79994 142980 79996
rect 142924 79942 142926 79994
rect 142926 79942 142978 79994
rect 142978 79942 142980 79994
rect 142924 79940 142980 79942
rect 142716 78426 142772 78428
rect 142716 78374 142718 78426
rect 142718 78374 142770 78426
rect 142770 78374 142772 78426
rect 142716 78372 142772 78374
rect 142820 78426 142876 78428
rect 142820 78374 142822 78426
rect 142822 78374 142874 78426
rect 142874 78374 142876 78426
rect 142820 78372 142876 78374
rect 142924 78426 142980 78428
rect 142924 78374 142926 78426
rect 142926 78374 142978 78426
rect 142978 78374 142980 78426
rect 142924 78372 142980 78374
rect 142716 76858 142772 76860
rect 142716 76806 142718 76858
rect 142718 76806 142770 76858
rect 142770 76806 142772 76858
rect 142716 76804 142772 76806
rect 142820 76858 142876 76860
rect 142820 76806 142822 76858
rect 142822 76806 142874 76858
rect 142874 76806 142876 76858
rect 142820 76804 142876 76806
rect 142924 76858 142980 76860
rect 142924 76806 142926 76858
rect 142926 76806 142978 76858
rect 142978 76806 142980 76858
rect 142924 76804 142980 76806
rect 142716 75290 142772 75292
rect 142716 75238 142718 75290
rect 142718 75238 142770 75290
rect 142770 75238 142772 75290
rect 142716 75236 142772 75238
rect 142820 75290 142876 75292
rect 142820 75238 142822 75290
rect 142822 75238 142874 75290
rect 142874 75238 142876 75290
rect 142820 75236 142876 75238
rect 142924 75290 142980 75292
rect 142924 75238 142926 75290
rect 142926 75238 142978 75290
rect 142978 75238 142980 75290
rect 142924 75236 142980 75238
rect 142716 73722 142772 73724
rect 142716 73670 142718 73722
rect 142718 73670 142770 73722
rect 142770 73670 142772 73722
rect 142716 73668 142772 73670
rect 142820 73722 142876 73724
rect 142820 73670 142822 73722
rect 142822 73670 142874 73722
rect 142874 73670 142876 73722
rect 142820 73668 142876 73670
rect 142924 73722 142980 73724
rect 142924 73670 142926 73722
rect 142926 73670 142978 73722
rect 142978 73670 142980 73722
rect 142924 73668 142980 73670
rect 142716 72154 142772 72156
rect 142716 72102 142718 72154
rect 142718 72102 142770 72154
rect 142770 72102 142772 72154
rect 142716 72100 142772 72102
rect 142820 72154 142876 72156
rect 142820 72102 142822 72154
rect 142822 72102 142874 72154
rect 142874 72102 142876 72154
rect 142820 72100 142876 72102
rect 142924 72154 142980 72156
rect 142924 72102 142926 72154
rect 142926 72102 142978 72154
rect 142978 72102 142980 72154
rect 142924 72100 142980 72102
rect 142716 70586 142772 70588
rect 142716 70534 142718 70586
rect 142718 70534 142770 70586
rect 142770 70534 142772 70586
rect 142716 70532 142772 70534
rect 142820 70586 142876 70588
rect 142820 70534 142822 70586
rect 142822 70534 142874 70586
rect 142874 70534 142876 70586
rect 142820 70532 142876 70534
rect 142924 70586 142980 70588
rect 142924 70534 142926 70586
rect 142926 70534 142978 70586
rect 142978 70534 142980 70586
rect 142924 70532 142980 70534
rect 142716 69018 142772 69020
rect 142716 68966 142718 69018
rect 142718 68966 142770 69018
rect 142770 68966 142772 69018
rect 142716 68964 142772 68966
rect 142820 69018 142876 69020
rect 142820 68966 142822 69018
rect 142822 68966 142874 69018
rect 142874 68966 142876 69018
rect 142820 68964 142876 68966
rect 142924 69018 142980 69020
rect 142924 68966 142926 69018
rect 142926 68966 142978 69018
rect 142978 68966 142980 69018
rect 142924 68964 142980 68966
rect 142716 67450 142772 67452
rect 142716 67398 142718 67450
rect 142718 67398 142770 67450
rect 142770 67398 142772 67450
rect 142716 67396 142772 67398
rect 142820 67450 142876 67452
rect 142820 67398 142822 67450
rect 142822 67398 142874 67450
rect 142874 67398 142876 67450
rect 142820 67396 142876 67398
rect 142924 67450 142980 67452
rect 142924 67398 142926 67450
rect 142926 67398 142978 67450
rect 142978 67398 142980 67450
rect 142924 67396 142980 67398
rect 142716 65882 142772 65884
rect 142716 65830 142718 65882
rect 142718 65830 142770 65882
rect 142770 65830 142772 65882
rect 142716 65828 142772 65830
rect 142820 65882 142876 65884
rect 142820 65830 142822 65882
rect 142822 65830 142874 65882
rect 142874 65830 142876 65882
rect 142820 65828 142876 65830
rect 142924 65882 142980 65884
rect 142924 65830 142926 65882
rect 142926 65830 142978 65882
rect 142978 65830 142980 65882
rect 142924 65828 142980 65830
rect 142716 64314 142772 64316
rect 142716 64262 142718 64314
rect 142718 64262 142770 64314
rect 142770 64262 142772 64314
rect 142716 64260 142772 64262
rect 142820 64314 142876 64316
rect 142820 64262 142822 64314
rect 142822 64262 142874 64314
rect 142874 64262 142876 64314
rect 142820 64260 142876 64262
rect 142924 64314 142980 64316
rect 142924 64262 142926 64314
rect 142926 64262 142978 64314
rect 142978 64262 142980 64314
rect 142924 64260 142980 64262
rect 142716 62746 142772 62748
rect 142716 62694 142718 62746
rect 142718 62694 142770 62746
rect 142770 62694 142772 62746
rect 142716 62692 142772 62694
rect 142820 62746 142876 62748
rect 142820 62694 142822 62746
rect 142822 62694 142874 62746
rect 142874 62694 142876 62746
rect 142820 62692 142876 62694
rect 142924 62746 142980 62748
rect 142924 62694 142926 62746
rect 142926 62694 142978 62746
rect 142978 62694 142980 62746
rect 142924 62692 142980 62694
rect 142716 61178 142772 61180
rect 142716 61126 142718 61178
rect 142718 61126 142770 61178
rect 142770 61126 142772 61178
rect 142716 61124 142772 61126
rect 142820 61178 142876 61180
rect 142820 61126 142822 61178
rect 142822 61126 142874 61178
rect 142874 61126 142876 61178
rect 142820 61124 142876 61126
rect 142924 61178 142980 61180
rect 142924 61126 142926 61178
rect 142926 61126 142978 61178
rect 142978 61126 142980 61178
rect 142924 61124 142980 61126
rect 142716 59610 142772 59612
rect 142716 59558 142718 59610
rect 142718 59558 142770 59610
rect 142770 59558 142772 59610
rect 142716 59556 142772 59558
rect 142820 59610 142876 59612
rect 142820 59558 142822 59610
rect 142822 59558 142874 59610
rect 142874 59558 142876 59610
rect 142820 59556 142876 59558
rect 142924 59610 142980 59612
rect 142924 59558 142926 59610
rect 142926 59558 142978 59610
rect 142978 59558 142980 59610
rect 142924 59556 142980 59558
rect 142716 58042 142772 58044
rect 142716 57990 142718 58042
rect 142718 57990 142770 58042
rect 142770 57990 142772 58042
rect 142716 57988 142772 57990
rect 142820 58042 142876 58044
rect 142820 57990 142822 58042
rect 142822 57990 142874 58042
rect 142874 57990 142876 58042
rect 142820 57988 142876 57990
rect 142924 58042 142980 58044
rect 142924 57990 142926 58042
rect 142926 57990 142978 58042
rect 142978 57990 142980 58042
rect 142924 57988 142980 57990
rect 142716 56474 142772 56476
rect 142716 56422 142718 56474
rect 142718 56422 142770 56474
rect 142770 56422 142772 56474
rect 142716 56420 142772 56422
rect 142820 56474 142876 56476
rect 142820 56422 142822 56474
rect 142822 56422 142874 56474
rect 142874 56422 142876 56474
rect 142820 56420 142876 56422
rect 142924 56474 142980 56476
rect 142924 56422 142926 56474
rect 142926 56422 142978 56474
rect 142978 56422 142980 56474
rect 142924 56420 142980 56422
rect 142716 54906 142772 54908
rect 142716 54854 142718 54906
rect 142718 54854 142770 54906
rect 142770 54854 142772 54906
rect 142716 54852 142772 54854
rect 142820 54906 142876 54908
rect 142820 54854 142822 54906
rect 142822 54854 142874 54906
rect 142874 54854 142876 54906
rect 142820 54852 142876 54854
rect 142924 54906 142980 54908
rect 142924 54854 142926 54906
rect 142926 54854 142978 54906
rect 142978 54854 142980 54906
rect 142924 54852 142980 54854
rect 142716 53338 142772 53340
rect 142716 53286 142718 53338
rect 142718 53286 142770 53338
rect 142770 53286 142772 53338
rect 142716 53284 142772 53286
rect 142820 53338 142876 53340
rect 142820 53286 142822 53338
rect 142822 53286 142874 53338
rect 142874 53286 142876 53338
rect 142820 53284 142876 53286
rect 142924 53338 142980 53340
rect 142924 53286 142926 53338
rect 142926 53286 142978 53338
rect 142978 53286 142980 53338
rect 142924 53284 142980 53286
rect 142716 51770 142772 51772
rect 142716 51718 142718 51770
rect 142718 51718 142770 51770
rect 142770 51718 142772 51770
rect 142716 51716 142772 51718
rect 142820 51770 142876 51772
rect 142820 51718 142822 51770
rect 142822 51718 142874 51770
rect 142874 51718 142876 51770
rect 142820 51716 142876 51718
rect 142924 51770 142980 51772
rect 142924 51718 142926 51770
rect 142926 51718 142978 51770
rect 142978 51718 142980 51770
rect 142924 51716 142980 51718
rect 142716 50202 142772 50204
rect 142716 50150 142718 50202
rect 142718 50150 142770 50202
rect 142770 50150 142772 50202
rect 142716 50148 142772 50150
rect 142820 50202 142876 50204
rect 142820 50150 142822 50202
rect 142822 50150 142874 50202
rect 142874 50150 142876 50202
rect 142820 50148 142876 50150
rect 142924 50202 142980 50204
rect 142924 50150 142926 50202
rect 142926 50150 142978 50202
rect 142978 50150 142980 50202
rect 142924 50148 142980 50150
rect 142716 48634 142772 48636
rect 142716 48582 142718 48634
rect 142718 48582 142770 48634
rect 142770 48582 142772 48634
rect 142716 48580 142772 48582
rect 142820 48634 142876 48636
rect 142820 48582 142822 48634
rect 142822 48582 142874 48634
rect 142874 48582 142876 48634
rect 142820 48580 142876 48582
rect 142924 48634 142980 48636
rect 142924 48582 142926 48634
rect 142926 48582 142978 48634
rect 142978 48582 142980 48634
rect 142924 48580 142980 48582
rect 142716 47066 142772 47068
rect 142716 47014 142718 47066
rect 142718 47014 142770 47066
rect 142770 47014 142772 47066
rect 142716 47012 142772 47014
rect 142820 47066 142876 47068
rect 142820 47014 142822 47066
rect 142822 47014 142874 47066
rect 142874 47014 142876 47066
rect 142820 47012 142876 47014
rect 142924 47066 142980 47068
rect 142924 47014 142926 47066
rect 142926 47014 142978 47066
rect 142978 47014 142980 47066
rect 142924 47012 142980 47014
rect 142716 45498 142772 45500
rect 142716 45446 142718 45498
rect 142718 45446 142770 45498
rect 142770 45446 142772 45498
rect 142716 45444 142772 45446
rect 142820 45498 142876 45500
rect 142820 45446 142822 45498
rect 142822 45446 142874 45498
rect 142874 45446 142876 45498
rect 142820 45444 142876 45446
rect 142924 45498 142980 45500
rect 142924 45446 142926 45498
rect 142926 45446 142978 45498
rect 142978 45446 142980 45498
rect 142924 45444 142980 45446
rect 142716 43930 142772 43932
rect 142716 43878 142718 43930
rect 142718 43878 142770 43930
rect 142770 43878 142772 43930
rect 142716 43876 142772 43878
rect 142820 43930 142876 43932
rect 142820 43878 142822 43930
rect 142822 43878 142874 43930
rect 142874 43878 142876 43930
rect 142820 43876 142876 43878
rect 142924 43930 142980 43932
rect 142924 43878 142926 43930
rect 142926 43878 142978 43930
rect 142978 43878 142980 43930
rect 142924 43876 142980 43878
rect 142716 42362 142772 42364
rect 142716 42310 142718 42362
rect 142718 42310 142770 42362
rect 142770 42310 142772 42362
rect 142716 42308 142772 42310
rect 142820 42362 142876 42364
rect 142820 42310 142822 42362
rect 142822 42310 142874 42362
rect 142874 42310 142876 42362
rect 142820 42308 142876 42310
rect 142924 42362 142980 42364
rect 142924 42310 142926 42362
rect 142926 42310 142978 42362
rect 142978 42310 142980 42362
rect 142924 42308 142980 42310
rect 142716 40794 142772 40796
rect 142716 40742 142718 40794
rect 142718 40742 142770 40794
rect 142770 40742 142772 40794
rect 142716 40740 142772 40742
rect 142820 40794 142876 40796
rect 142820 40742 142822 40794
rect 142822 40742 142874 40794
rect 142874 40742 142876 40794
rect 142820 40740 142876 40742
rect 142924 40794 142980 40796
rect 142924 40742 142926 40794
rect 142926 40742 142978 40794
rect 142978 40742 142980 40794
rect 142924 40740 142980 40742
rect 142716 39226 142772 39228
rect 142716 39174 142718 39226
rect 142718 39174 142770 39226
rect 142770 39174 142772 39226
rect 142716 39172 142772 39174
rect 142820 39226 142876 39228
rect 142820 39174 142822 39226
rect 142822 39174 142874 39226
rect 142874 39174 142876 39226
rect 142820 39172 142876 39174
rect 142924 39226 142980 39228
rect 142924 39174 142926 39226
rect 142926 39174 142978 39226
rect 142978 39174 142980 39226
rect 142924 39172 142980 39174
rect 142716 37658 142772 37660
rect 142716 37606 142718 37658
rect 142718 37606 142770 37658
rect 142770 37606 142772 37658
rect 142716 37604 142772 37606
rect 142820 37658 142876 37660
rect 142820 37606 142822 37658
rect 142822 37606 142874 37658
rect 142874 37606 142876 37658
rect 142820 37604 142876 37606
rect 142924 37658 142980 37660
rect 142924 37606 142926 37658
rect 142926 37606 142978 37658
rect 142978 37606 142980 37658
rect 142924 37604 142980 37606
rect 142716 36090 142772 36092
rect 142716 36038 142718 36090
rect 142718 36038 142770 36090
rect 142770 36038 142772 36090
rect 142716 36036 142772 36038
rect 142820 36090 142876 36092
rect 142820 36038 142822 36090
rect 142822 36038 142874 36090
rect 142874 36038 142876 36090
rect 142820 36036 142876 36038
rect 142924 36090 142980 36092
rect 142924 36038 142926 36090
rect 142926 36038 142978 36090
rect 142978 36038 142980 36090
rect 142924 36036 142980 36038
rect 142716 34522 142772 34524
rect 142716 34470 142718 34522
rect 142718 34470 142770 34522
rect 142770 34470 142772 34522
rect 142716 34468 142772 34470
rect 142820 34522 142876 34524
rect 142820 34470 142822 34522
rect 142822 34470 142874 34522
rect 142874 34470 142876 34522
rect 142820 34468 142876 34470
rect 142924 34522 142980 34524
rect 142924 34470 142926 34522
rect 142926 34470 142978 34522
rect 142978 34470 142980 34522
rect 142924 34468 142980 34470
rect 142716 32954 142772 32956
rect 142716 32902 142718 32954
rect 142718 32902 142770 32954
rect 142770 32902 142772 32954
rect 142716 32900 142772 32902
rect 142820 32954 142876 32956
rect 142820 32902 142822 32954
rect 142822 32902 142874 32954
rect 142874 32902 142876 32954
rect 142820 32900 142876 32902
rect 142924 32954 142980 32956
rect 142924 32902 142926 32954
rect 142926 32902 142978 32954
rect 142978 32902 142980 32954
rect 142924 32900 142980 32902
rect 142716 31386 142772 31388
rect 142716 31334 142718 31386
rect 142718 31334 142770 31386
rect 142770 31334 142772 31386
rect 142716 31332 142772 31334
rect 142820 31386 142876 31388
rect 142820 31334 142822 31386
rect 142822 31334 142874 31386
rect 142874 31334 142876 31386
rect 142820 31332 142876 31334
rect 142924 31386 142980 31388
rect 142924 31334 142926 31386
rect 142926 31334 142978 31386
rect 142978 31334 142980 31386
rect 142924 31332 142980 31334
rect 142716 29818 142772 29820
rect 142716 29766 142718 29818
rect 142718 29766 142770 29818
rect 142770 29766 142772 29818
rect 142716 29764 142772 29766
rect 142820 29818 142876 29820
rect 142820 29766 142822 29818
rect 142822 29766 142874 29818
rect 142874 29766 142876 29818
rect 142820 29764 142876 29766
rect 142924 29818 142980 29820
rect 142924 29766 142926 29818
rect 142926 29766 142978 29818
rect 142978 29766 142980 29818
rect 142924 29764 142980 29766
rect 142716 28250 142772 28252
rect 142716 28198 142718 28250
rect 142718 28198 142770 28250
rect 142770 28198 142772 28250
rect 142716 28196 142772 28198
rect 142820 28250 142876 28252
rect 142820 28198 142822 28250
rect 142822 28198 142874 28250
rect 142874 28198 142876 28250
rect 142820 28196 142876 28198
rect 142924 28250 142980 28252
rect 142924 28198 142926 28250
rect 142926 28198 142978 28250
rect 142978 28198 142980 28250
rect 142924 28196 142980 28198
rect 142716 26682 142772 26684
rect 142716 26630 142718 26682
rect 142718 26630 142770 26682
rect 142770 26630 142772 26682
rect 142716 26628 142772 26630
rect 142820 26682 142876 26684
rect 142820 26630 142822 26682
rect 142822 26630 142874 26682
rect 142874 26630 142876 26682
rect 142820 26628 142876 26630
rect 142924 26682 142980 26684
rect 142924 26630 142926 26682
rect 142926 26630 142978 26682
rect 142978 26630 142980 26682
rect 142924 26628 142980 26630
rect 142716 25114 142772 25116
rect 142716 25062 142718 25114
rect 142718 25062 142770 25114
rect 142770 25062 142772 25114
rect 142716 25060 142772 25062
rect 142820 25114 142876 25116
rect 142820 25062 142822 25114
rect 142822 25062 142874 25114
rect 142874 25062 142876 25114
rect 142820 25060 142876 25062
rect 142924 25114 142980 25116
rect 142924 25062 142926 25114
rect 142926 25062 142978 25114
rect 142978 25062 142980 25114
rect 142924 25060 142980 25062
rect 142716 23546 142772 23548
rect 142716 23494 142718 23546
rect 142718 23494 142770 23546
rect 142770 23494 142772 23546
rect 142716 23492 142772 23494
rect 142820 23546 142876 23548
rect 142820 23494 142822 23546
rect 142822 23494 142874 23546
rect 142874 23494 142876 23546
rect 142820 23492 142876 23494
rect 142924 23546 142980 23548
rect 142924 23494 142926 23546
rect 142926 23494 142978 23546
rect 142978 23494 142980 23546
rect 142924 23492 142980 23494
rect 142716 21978 142772 21980
rect 142716 21926 142718 21978
rect 142718 21926 142770 21978
rect 142770 21926 142772 21978
rect 142716 21924 142772 21926
rect 142820 21978 142876 21980
rect 142820 21926 142822 21978
rect 142822 21926 142874 21978
rect 142874 21926 142876 21978
rect 142820 21924 142876 21926
rect 142924 21978 142980 21980
rect 142924 21926 142926 21978
rect 142926 21926 142978 21978
rect 142978 21926 142980 21978
rect 142924 21924 142980 21926
rect 142716 20410 142772 20412
rect 142716 20358 142718 20410
rect 142718 20358 142770 20410
rect 142770 20358 142772 20410
rect 142716 20356 142772 20358
rect 142820 20410 142876 20412
rect 142820 20358 142822 20410
rect 142822 20358 142874 20410
rect 142874 20358 142876 20410
rect 142820 20356 142876 20358
rect 142924 20410 142980 20412
rect 142924 20358 142926 20410
rect 142926 20358 142978 20410
rect 142978 20358 142980 20410
rect 142924 20356 142980 20358
rect 140700 19292 140756 19348
rect 142716 18842 142772 18844
rect 142716 18790 142718 18842
rect 142718 18790 142770 18842
rect 142770 18790 142772 18842
rect 142716 18788 142772 18790
rect 142820 18842 142876 18844
rect 142820 18790 142822 18842
rect 142822 18790 142874 18842
rect 142874 18790 142876 18842
rect 142820 18788 142876 18790
rect 142924 18842 142980 18844
rect 142924 18790 142926 18842
rect 142926 18790 142978 18842
rect 142978 18790 142980 18842
rect 142924 18788 142980 18790
rect 136892 17612 136948 17668
rect 137228 17836 137284 17892
rect 136780 8540 136836 8596
rect 137116 13916 137172 13972
rect 136668 8204 136724 8260
rect 135884 6690 135940 6692
rect 135884 6638 135886 6690
rect 135886 6638 135938 6690
rect 135938 6638 135940 6690
rect 135884 6636 135940 6638
rect 135772 6412 135828 6468
rect 135772 6018 135828 6020
rect 135772 5966 135774 6018
rect 135774 5966 135826 6018
rect 135826 5966 135828 6018
rect 135772 5964 135828 5966
rect 135548 5404 135604 5460
rect 135436 5292 135492 5348
rect 136220 6188 136276 6244
rect 135996 5852 136052 5908
rect 135660 5010 135716 5012
rect 135660 4958 135662 5010
rect 135662 4958 135714 5010
rect 135714 4958 135716 5010
rect 135660 4956 135716 4958
rect 135324 4732 135380 4788
rect 135660 4508 135716 4564
rect 135212 3612 135268 3668
rect 135436 3612 135492 3668
rect 135324 3500 135380 3556
rect 134092 3052 134148 3108
rect 134092 2492 134148 2548
rect 136108 5068 136164 5124
rect 135884 4732 135940 4788
rect 135772 3052 135828 3108
rect 135884 4508 135940 4564
rect 136108 4450 136164 4452
rect 136108 4398 136110 4450
rect 136110 4398 136162 4450
rect 136162 4398 136164 4450
rect 136108 4396 136164 4398
rect 135996 2380 136052 2436
rect 136220 3724 136276 3780
rect 136332 3836 136388 3892
rect 136332 3442 136388 3444
rect 136332 3390 136334 3442
rect 136334 3390 136386 3442
rect 136386 3390 136388 3442
rect 136332 3388 136388 3390
rect 136108 1596 136164 1652
rect 136668 5740 136724 5796
rect 136668 4956 136724 5012
rect 136892 6636 136948 6692
rect 137004 6130 137060 6132
rect 137004 6078 137006 6130
rect 137006 6078 137058 6130
rect 137058 6078 137060 6130
rect 137004 6076 137060 6078
rect 136780 4620 136836 4676
rect 142716 17274 142772 17276
rect 142716 17222 142718 17274
rect 142718 17222 142770 17274
rect 142770 17222 142772 17274
rect 142716 17220 142772 17222
rect 142820 17274 142876 17276
rect 142820 17222 142822 17274
rect 142822 17222 142874 17274
rect 142874 17222 142876 17274
rect 142820 17220 142876 17222
rect 142924 17274 142980 17276
rect 142924 17222 142926 17274
rect 142926 17222 142978 17274
rect 142978 17222 142980 17274
rect 142924 17220 142980 17222
rect 142716 15706 142772 15708
rect 142716 15654 142718 15706
rect 142718 15654 142770 15706
rect 142770 15654 142772 15706
rect 142716 15652 142772 15654
rect 142820 15706 142876 15708
rect 142820 15654 142822 15706
rect 142822 15654 142874 15706
rect 142874 15654 142876 15706
rect 142820 15652 142876 15654
rect 142924 15706 142980 15708
rect 142924 15654 142926 15706
rect 142926 15654 142978 15706
rect 142978 15654 142980 15706
rect 142924 15652 142980 15654
rect 142604 15372 142660 15428
rect 141820 13804 141876 13860
rect 141372 13692 141428 13748
rect 139132 8876 139188 8932
rect 137788 8540 137844 8596
rect 137340 6972 137396 7028
rect 137452 7308 137508 7364
rect 137340 6636 137396 6692
rect 137228 6466 137284 6468
rect 137228 6414 137230 6466
rect 137230 6414 137282 6466
rect 137282 6414 137284 6466
rect 137228 6412 137284 6414
rect 137340 5404 137396 5460
rect 137340 5010 137396 5012
rect 137340 4958 137342 5010
rect 137342 4958 137394 5010
rect 137394 4958 137396 5010
rect 137340 4956 137396 4958
rect 138908 8092 138964 8148
rect 138012 7756 138068 7812
rect 137564 6748 137620 6804
rect 137564 5404 137620 5460
rect 137676 6188 137732 6244
rect 137788 5794 137844 5796
rect 137788 5742 137790 5794
rect 137790 5742 137842 5794
rect 137842 5742 137844 5794
rect 137788 5740 137844 5742
rect 137676 5292 137732 5348
rect 137788 5234 137844 5236
rect 137788 5182 137790 5234
rect 137790 5182 137842 5234
rect 137842 5182 137844 5234
rect 137788 5180 137844 5182
rect 137900 5010 137956 5012
rect 137900 4958 137902 5010
rect 137902 4958 137954 5010
rect 137954 4958 137956 5010
rect 137900 4956 137956 4958
rect 138796 7308 138852 7364
rect 138236 7084 138292 7140
rect 138236 6748 138292 6804
rect 138124 5852 138180 5908
rect 138684 6636 138740 6692
rect 138684 6076 138740 6132
rect 138348 5010 138404 5012
rect 138348 4958 138350 5010
rect 138350 4958 138402 5010
rect 138402 4958 138404 5010
rect 138348 4956 138404 4958
rect 137116 4226 137172 4228
rect 137116 4174 137118 4226
rect 137118 4174 137170 4226
rect 137170 4174 137172 4226
rect 137116 4172 137172 4174
rect 137340 3948 137396 4004
rect 137116 3724 137172 3780
rect 137340 3724 137396 3780
rect 137788 3948 137844 4004
rect 137004 3388 137060 3444
rect 136892 3330 136948 3332
rect 136892 3278 136894 3330
rect 136894 3278 136946 3330
rect 136946 3278 136948 3330
rect 136892 3276 136948 3278
rect 136668 2604 136724 2660
rect 138012 3724 138068 3780
rect 138572 4508 138628 4564
rect 138796 4844 138852 4900
rect 138684 4284 138740 4340
rect 138572 4114 138628 4116
rect 138572 4062 138574 4114
rect 138574 4062 138626 4114
rect 138626 4062 138628 4114
rect 138572 4060 138628 4062
rect 137676 924 137732 980
rect 138908 3836 138964 3892
rect 140476 8764 140532 8820
rect 139132 6578 139188 6580
rect 139132 6526 139134 6578
rect 139134 6526 139186 6578
rect 139186 6526 139188 6578
rect 139132 6524 139188 6526
rect 139132 6188 139188 6244
rect 139356 6412 139412 6468
rect 139132 4844 139188 4900
rect 139020 3724 139076 3780
rect 139132 3388 139188 3444
rect 139804 6524 139860 6580
rect 140140 6524 140196 6580
rect 140028 6188 140084 6244
rect 139804 5682 139860 5684
rect 139804 5630 139806 5682
rect 139806 5630 139858 5682
rect 139858 5630 139860 5682
rect 139804 5628 139860 5630
rect 139692 4620 139748 4676
rect 139468 4172 139524 4228
rect 139692 4172 139748 4228
rect 139244 2828 139300 2884
rect 139916 3500 139972 3556
rect 139916 3052 139972 3108
rect 140476 7362 140532 7364
rect 140476 7310 140478 7362
rect 140478 7310 140530 7362
rect 140530 7310 140532 7362
rect 140476 7308 140532 7310
rect 140924 6300 140980 6356
rect 140700 6188 140756 6244
rect 140812 6130 140868 6132
rect 140812 6078 140814 6130
rect 140814 6078 140866 6130
rect 140866 6078 140868 6130
rect 140812 6076 140868 6078
rect 140588 5628 140644 5684
rect 140924 5740 140980 5796
rect 140924 4620 140980 4676
rect 140252 4284 140308 4340
rect 140252 3554 140308 3556
rect 140252 3502 140254 3554
rect 140254 3502 140306 3554
rect 140306 3502 140308 3554
rect 140252 3500 140308 3502
rect 140588 4338 140644 4340
rect 140588 4286 140590 4338
rect 140590 4286 140642 4338
rect 140642 4286 140644 4338
rect 140588 4284 140644 4286
rect 140364 3276 140420 3332
rect 140476 3724 140532 3780
rect 140140 3164 140196 3220
rect 139692 2380 139748 2436
rect 140700 812 140756 868
rect 141260 6748 141316 6804
rect 141260 5010 141316 5012
rect 141260 4958 141262 5010
rect 141262 4958 141314 5010
rect 141314 4958 141316 5010
rect 141260 4956 141316 4958
rect 141708 6188 141764 6244
rect 142492 12348 142548 12404
rect 141148 3948 141204 4004
rect 141596 4732 141652 4788
rect 141708 4562 141764 4564
rect 141708 4510 141710 4562
rect 141710 4510 141762 4562
rect 141762 4510 141764 4562
rect 141708 4508 141764 4510
rect 141820 4338 141876 4340
rect 141820 4286 141822 4338
rect 141822 4286 141874 4338
rect 141874 4286 141876 4338
rect 141820 4284 141876 4286
rect 142044 6636 142100 6692
rect 142044 5068 142100 5124
rect 142268 6300 142324 6356
rect 142380 6412 142436 6468
rect 142716 14138 142772 14140
rect 142716 14086 142718 14138
rect 142718 14086 142770 14138
rect 142770 14086 142772 14138
rect 142716 14084 142772 14086
rect 142820 14138 142876 14140
rect 142820 14086 142822 14138
rect 142822 14086 142874 14138
rect 142874 14086 142876 14138
rect 142820 14084 142876 14086
rect 142924 14138 142980 14140
rect 142924 14086 142926 14138
rect 142926 14086 142978 14138
rect 142978 14086 142980 14138
rect 142924 14084 142980 14086
rect 143724 12908 143780 12964
rect 142716 12570 142772 12572
rect 142716 12518 142718 12570
rect 142718 12518 142770 12570
rect 142770 12518 142772 12570
rect 142716 12516 142772 12518
rect 142820 12570 142876 12572
rect 142820 12518 142822 12570
rect 142822 12518 142874 12570
rect 142874 12518 142876 12570
rect 142820 12516 142876 12518
rect 142924 12570 142980 12572
rect 142924 12518 142926 12570
rect 142926 12518 142978 12570
rect 142978 12518 142980 12570
rect 142924 12516 142980 12518
rect 142716 11002 142772 11004
rect 142716 10950 142718 11002
rect 142718 10950 142770 11002
rect 142770 10950 142772 11002
rect 142716 10948 142772 10950
rect 142820 11002 142876 11004
rect 142820 10950 142822 11002
rect 142822 10950 142874 11002
rect 142874 10950 142876 11002
rect 142820 10948 142876 10950
rect 142924 11002 142980 11004
rect 142924 10950 142926 11002
rect 142926 10950 142978 11002
rect 142978 10950 142980 11002
rect 142924 10948 142980 10950
rect 142716 9434 142772 9436
rect 142716 9382 142718 9434
rect 142718 9382 142770 9434
rect 142770 9382 142772 9434
rect 142716 9380 142772 9382
rect 142820 9434 142876 9436
rect 142820 9382 142822 9434
rect 142822 9382 142874 9434
rect 142874 9382 142876 9434
rect 142820 9380 142876 9382
rect 142924 9434 142980 9436
rect 142924 9382 142926 9434
rect 142926 9382 142978 9434
rect 142978 9382 142980 9434
rect 142924 9380 142980 9382
rect 142716 7866 142772 7868
rect 142716 7814 142718 7866
rect 142718 7814 142770 7866
rect 142770 7814 142772 7866
rect 142716 7812 142772 7814
rect 142820 7866 142876 7868
rect 142820 7814 142822 7866
rect 142822 7814 142874 7866
rect 142874 7814 142876 7866
rect 142820 7812 142876 7814
rect 142924 7866 142980 7868
rect 142924 7814 142926 7866
rect 142926 7814 142978 7866
rect 142978 7814 142980 7866
rect 142924 7812 142980 7814
rect 142716 6636 142772 6692
rect 142604 6466 142660 6468
rect 142604 6414 142606 6466
rect 142606 6414 142658 6466
rect 142658 6414 142660 6466
rect 142604 6412 142660 6414
rect 143052 6466 143108 6468
rect 143052 6414 143054 6466
rect 143054 6414 143106 6466
rect 143106 6414 143108 6466
rect 143052 6412 143108 6414
rect 142716 6298 142772 6300
rect 142716 6246 142718 6298
rect 142718 6246 142770 6298
rect 142770 6246 142772 6298
rect 142716 6244 142772 6246
rect 142820 6298 142876 6300
rect 142820 6246 142822 6298
rect 142822 6246 142874 6298
rect 142874 6246 142876 6298
rect 142820 6244 142876 6246
rect 142924 6298 142980 6300
rect 142924 6246 142926 6298
rect 142926 6246 142978 6298
rect 142978 6246 142980 6298
rect 142924 6244 142980 6246
rect 142380 6018 142436 6020
rect 142380 5966 142382 6018
rect 142382 5966 142434 6018
rect 142434 5966 142436 6018
rect 142380 5964 142436 5966
rect 142268 5180 142324 5236
rect 142716 5628 142772 5684
rect 142156 4620 142212 4676
rect 142716 4730 142772 4732
rect 142716 4678 142718 4730
rect 142718 4678 142770 4730
rect 142770 4678 142772 4730
rect 142716 4676 142772 4678
rect 142820 4730 142876 4732
rect 142820 4678 142822 4730
rect 142822 4678 142874 4730
rect 142874 4678 142876 4730
rect 142820 4676 142876 4678
rect 142924 4730 142980 4732
rect 142924 4678 142926 4730
rect 142926 4678 142978 4730
rect 142978 4678 142980 4730
rect 142924 4676 142980 4678
rect 143052 4508 143108 4564
rect 142268 4226 142324 4228
rect 142268 4174 142270 4226
rect 142270 4174 142322 4226
rect 142322 4174 142324 4226
rect 142268 4172 142324 4174
rect 143052 4226 143108 4228
rect 143052 4174 143054 4226
rect 143054 4174 143106 4226
rect 143106 4174 143108 4226
rect 143052 4172 143108 4174
rect 142604 3612 142660 3668
rect 142156 3500 142212 3556
rect 142044 3442 142100 3444
rect 142044 3390 142046 3442
rect 142046 3390 142098 3442
rect 142098 3390 142100 3442
rect 142044 3388 142100 3390
rect 141036 2828 141092 2884
rect 142940 3330 142996 3332
rect 142940 3278 142942 3330
rect 142942 3278 142994 3330
rect 142994 3278 142996 3330
rect 142940 3276 142996 3278
rect 142716 3162 142772 3164
rect 142716 3110 142718 3162
rect 142718 3110 142770 3162
rect 142770 3110 142772 3162
rect 142716 3108 142772 3110
rect 142820 3162 142876 3164
rect 142820 3110 142822 3162
rect 142822 3110 142874 3162
rect 142874 3110 142876 3162
rect 142820 3108 142876 3110
rect 142924 3162 142980 3164
rect 142924 3110 142926 3162
rect 142926 3110 142978 3162
rect 142978 3110 142980 3162
rect 142924 3108 142980 3110
rect 143388 5740 143444 5796
rect 143276 4620 143332 4676
rect 143276 3724 143332 3780
rect 143500 4172 143556 4228
rect 145964 12124 146020 12180
rect 143948 7644 144004 7700
rect 143724 5740 143780 5796
rect 143724 5516 143780 5572
rect 143724 4732 143780 4788
rect 143724 4172 143780 4228
rect 143948 5628 144004 5684
rect 144060 5516 144116 5572
rect 144508 5964 144564 6020
rect 143948 5346 144004 5348
rect 143948 5294 143950 5346
rect 143950 5294 144002 5346
rect 144002 5294 144004 5346
rect 143948 5292 144004 5294
rect 144508 5292 144564 5348
rect 144060 5122 144116 5124
rect 144060 5070 144062 5122
rect 144062 5070 144114 5122
rect 144114 5070 144116 5122
rect 144060 5068 144116 5070
rect 143836 3724 143892 3780
rect 143612 3500 143668 3556
rect 143388 1036 143444 1092
rect 143724 3388 143780 3444
rect 144060 4562 144116 4564
rect 144060 4510 144062 4562
rect 144062 4510 144114 4562
rect 144114 4510 144116 4562
rect 144060 4508 144116 4510
rect 144284 3948 144340 4004
rect 144172 3554 144228 3556
rect 144172 3502 144174 3554
rect 144174 3502 144226 3554
rect 144226 3502 144228 3554
rect 144172 3500 144228 3502
rect 143948 3276 144004 3332
rect 143836 2828 143892 2884
rect 145180 6860 145236 6916
rect 144732 3612 144788 3668
rect 144956 6076 145012 6132
rect 145292 6018 145348 6020
rect 145292 5966 145294 6018
rect 145294 5966 145346 6018
rect 145346 5966 145348 6018
rect 145292 5964 145348 5966
rect 145180 5740 145236 5796
rect 145292 5010 145348 5012
rect 145292 4958 145294 5010
rect 145294 4958 145346 5010
rect 145346 4958 145348 5010
rect 145292 4956 145348 4958
rect 145180 4620 145236 4676
rect 145068 4338 145124 4340
rect 145068 4286 145070 4338
rect 145070 4286 145122 4338
rect 145122 4286 145124 4338
rect 145068 4284 145124 4286
rect 145740 6466 145796 6468
rect 145740 6414 145742 6466
rect 145742 6414 145794 6466
rect 145794 6414 145796 6466
rect 145740 6412 145796 6414
rect 145740 5964 145796 6020
rect 145516 4956 145572 5012
rect 145180 3724 145236 3780
rect 144956 3612 145012 3668
rect 145852 4732 145908 4788
rect 154700 116450 154756 116452
rect 154700 116398 154702 116450
rect 154702 116398 154754 116450
rect 154754 116398 154756 116450
rect 154700 116396 154756 116398
rect 155372 116956 155428 117012
rect 158076 116842 158132 116844
rect 158076 116790 158078 116842
rect 158078 116790 158130 116842
rect 158130 116790 158132 116842
rect 158076 116788 158132 116790
rect 158180 116842 158236 116844
rect 158180 116790 158182 116842
rect 158182 116790 158234 116842
rect 158234 116790 158236 116842
rect 158180 116788 158236 116790
rect 158284 116842 158340 116844
rect 158284 116790 158286 116842
rect 158286 116790 158338 116842
rect 158338 116790 158340 116842
rect 158284 116788 158340 116790
rect 162876 116620 162932 116676
rect 163772 116620 163828 116676
rect 167580 117068 167636 117124
rect 168476 117068 168532 117124
rect 164444 116284 164500 116340
rect 164892 116338 164948 116340
rect 164892 116286 164894 116338
rect 164894 116286 164946 116338
rect 164946 116286 164948 116338
rect 164892 116284 164948 116286
rect 172284 116620 172340 116676
rect 173068 116620 173124 116676
rect 170940 116396 170996 116452
rect 169148 116284 169204 116340
rect 170380 116338 170436 116340
rect 170380 116286 170382 116338
rect 170382 116286 170434 116338
rect 170434 116286 170436 116338
rect 170380 116284 170436 116286
rect 172284 116450 172340 116452
rect 172284 116398 172286 116450
rect 172286 116398 172338 116450
rect 172338 116398 172340 116450
rect 172284 116396 172340 116398
rect 173436 116058 173492 116060
rect 173436 116006 173438 116058
rect 173438 116006 173490 116058
rect 173490 116006 173492 116058
rect 173436 116004 173492 116006
rect 173540 116058 173596 116060
rect 173540 116006 173542 116058
rect 173542 116006 173594 116058
rect 173594 116006 173596 116058
rect 173540 116004 173596 116006
rect 173644 116058 173700 116060
rect 173644 116006 173646 116058
rect 173646 116006 173698 116058
rect 173698 116006 173700 116058
rect 173644 116004 173700 116006
rect 178108 115890 178164 115892
rect 178108 115838 178110 115890
rect 178110 115838 178162 115890
rect 178162 115838 178164 115890
rect 178108 115836 178164 115838
rect 178556 115836 178612 115892
rect 152124 115666 152180 115668
rect 152124 115614 152126 115666
rect 152126 115614 152178 115666
rect 152178 115614 152180 115666
rect 152124 115612 152180 115614
rect 153244 115666 153300 115668
rect 153244 115614 153246 115666
rect 153246 115614 153298 115666
rect 153298 115614 153300 115666
rect 153244 115612 153300 115614
rect 157276 115666 157332 115668
rect 157276 115614 157278 115666
rect 157278 115614 157330 115666
rect 157330 115614 157332 115666
rect 157276 115612 157332 115614
rect 157836 115666 157892 115668
rect 157836 115614 157838 115666
rect 157838 115614 157890 115666
rect 157890 115614 157892 115666
rect 157836 115612 157892 115614
rect 161980 115666 162036 115668
rect 161980 115614 161982 115666
rect 161982 115614 162034 115666
rect 162034 115614 162036 115666
rect 161980 115612 162036 115614
rect 162540 115666 162596 115668
rect 162540 115614 162542 115666
rect 162542 115614 162594 115666
rect 162594 115614 162596 115666
rect 162540 115612 162596 115614
rect 166684 115666 166740 115668
rect 166684 115614 166686 115666
rect 166686 115614 166738 115666
rect 166738 115614 166740 115666
rect 166684 115612 166740 115614
rect 167244 115666 167300 115668
rect 167244 115614 167246 115666
rect 167246 115614 167298 115666
rect 167298 115614 167300 115666
rect 167244 115612 167300 115614
rect 170044 115666 170100 115668
rect 170044 115614 170046 115666
rect 170046 115614 170098 115666
rect 170098 115614 170100 115666
rect 170044 115612 170100 115614
rect 170604 115666 170660 115668
rect 170604 115614 170606 115666
rect 170606 115614 170658 115666
rect 170658 115614 170660 115666
rect 170604 115612 170660 115614
rect 158076 115274 158132 115276
rect 158076 115222 158078 115274
rect 158078 115222 158130 115274
rect 158130 115222 158132 115274
rect 158076 115220 158132 115222
rect 158180 115274 158236 115276
rect 158180 115222 158182 115274
rect 158182 115222 158234 115274
rect 158234 115222 158236 115274
rect 158180 115220 158236 115222
rect 158284 115274 158340 115276
rect 158284 115222 158286 115274
rect 158286 115222 158338 115274
rect 158338 115222 158340 115274
rect 158284 115220 158340 115222
rect 173436 114490 173492 114492
rect 173436 114438 173438 114490
rect 173438 114438 173490 114490
rect 173490 114438 173492 114490
rect 173436 114436 173492 114438
rect 173540 114490 173596 114492
rect 173540 114438 173542 114490
rect 173542 114438 173594 114490
rect 173594 114438 173596 114490
rect 173540 114436 173596 114438
rect 173644 114490 173700 114492
rect 173644 114438 173646 114490
rect 173646 114438 173698 114490
rect 173698 114438 173700 114490
rect 173644 114436 173700 114438
rect 158076 113706 158132 113708
rect 158076 113654 158078 113706
rect 158078 113654 158130 113706
rect 158130 113654 158132 113706
rect 158076 113652 158132 113654
rect 158180 113706 158236 113708
rect 158180 113654 158182 113706
rect 158182 113654 158234 113706
rect 158234 113654 158236 113706
rect 158180 113652 158236 113654
rect 158284 113706 158340 113708
rect 158284 113654 158286 113706
rect 158286 113654 158338 113706
rect 158338 113654 158340 113706
rect 158284 113652 158340 113654
rect 173436 112922 173492 112924
rect 173436 112870 173438 112922
rect 173438 112870 173490 112922
rect 173490 112870 173492 112922
rect 173436 112868 173492 112870
rect 173540 112922 173596 112924
rect 173540 112870 173542 112922
rect 173542 112870 173594 112922
rect 173594 112870 173596 112922
rect 173540 112868 173596 112870
rect 173644 112922 173700 112924
rect 173644 112870 173646 112922
rect 173646 112870 173698 112922
rect 173698 112870 173700 112922
rect 173644 112868 173700 112870
rect 158076 112138 158132 112140
rect 158076 112086 158078 112138
rect 158078 112086 158130 112138
rect 158130 112086 158132 112138
rect 158076 112084 158132 112086
rect 158180 112138 158236 112140
rect 158180 112086 158182 112138
rect 158182 112086 158234 112138
rect 158234 112086 158236 112138
rect 158180 112084 158236 112086
rect 158284 112138 158340 112140
rect 158284 112086 158286 112138
rect 158286 112086 158338 112138
rect 158338 112086 158340 112138
rect 158284 112084 158340 112086
rect 173436 111354 173492 111356
rect 173436 111302 173438 111354
rect 173438 111302 173490 111354
rect 173490 111302 173492 111354
rect 173436 111300 173492 111302
rect 173540 111354 173596 111356
rect 173540 111302 173542 111354
rect 173542 111302 173594 111354
rect 173594 111302 173596 111354
rect 173540 111300 173596 111302
rect 173644 111354 173700 111356
rect 173644 111302 173646 111354
rect 173646 111302 173698 111354
rect 173698 111302 173700 111354
rect 173644 111300 173700 111302
rect 158076 110570 158132 110572
rect 158076 110518 158078 110570
rect 158078 110518 158130 110570
rect 158130 110518 158132 110570
rect 158076 110516 158132 110518
rect 158180 110570 158236 110572
rect 158180 110518 158182 110570
rect 158182 110518 158234 110570
rect 158234 110518 158236 110570
rect 158180 110516 158236 110518
rect 158284 110570 158340 110572
rect 158284 110518 158286 110570
rect 158286 110518 158338 110570
rect 158338 110518 158340 110570
rect 158284 110516 158340 110518
rect 173436 109786 173492 109788
rect 173436 109734 173438 109786
rect 173438 109734 173490 109786
rect 173490 109734 173492 109786
rect 173436 109732 173492 109734
rect 173540 109786 173596 109788
rect 173540 109734 173542 109786
rect 173542 109734 173594 109786
rect 173594 109734 173596 109786
rect 173540 109732 173596 109734
rect 173644 109786 173700 109788
rect 173644 109734 173646 109786
rect 173646 109734 173698 109786
rect 173698 109734 173700 109786
rect 173644 109732 173700 109734
rect 158076 109002 158132 109004
rect 158076 108950 158078 109002
rect 158078 108950 158130 109002
rect 158130 108950 158132 109002
rect 158076 108948 158132 108950
rect 158180 109002 158236 109004
rect 158180 108950 158182 109002
rect 158182 108950 158234 109002
rect 158234 108950 158236 109002
rect 158180 108948 158236 108950
rect 158284 109002 158340 109004
rect 158284 108950 158286 109002
rect 158286 108950 158338 109002
rect 158338 108950 158340 109002
rect 158284 108948 158340 108950
rect 173436 108218 173492 108220
rect 173436 108166 173438 108218
rect 173438 108166 173490 108218
rect 173490 108166 173492 108218
rect 173436 108164 173492 108166
rect 173540 108218 173596 108220
rect 173540 108166 173542 108218
rect 173542 108166 173594 108218
rect 173594 108166 173596 108218
rect 173540 108164 173596 108166
rect 173644 108218 173700 108220
rect 173644 108166 173646 108218
rect 173646 108166 173698 108218
rect 173698 108166 173700 108218
rect 173644 108164 173700 108166
rect 158076 107434 158132 107436
rect 158076 107382 158078 107434
rect 158078 107382 158130 107434
rect 158130 107382 158132 107434
rect 158076 107380 158132 107382
rect 158180 107434 158236 107436
rect 158180 107382 158182 107434
rect 158182 107382 158234 107434
rect 158234 107382 158236 107434
rect 158180 107380 158236 107382
rect 158284 107434 158340 107436
rect 158284 107382 158286 107434
rect 158286 107382 158338 107434
rect 158338 107382 158340 107434
rect 158284 107380 158340 107382
rect 173436 106650 173492 106652
rect 173436 106598 173438 106650
rect 173438 106598 173490 106650
rect 173490 106598 173492 106650
rect 173436 106596 173492 106598
rect 173540 106650 173596 106652
rect 173540 106598 173542 106650
rect 173542 106598 173594 106650
rect 173594 106598 173596 106650
rect 173540 106596 173596 106598
rect 173644 106650 173700 106652
rect 173644 106598 173646 106650
rect 173646 106598 173698 106650
rect 173698 106598 173700 106650
rect 173644 106596 173700 106598
rect 158076 105866 158132 105868
rect 158076 105814 158078 105866
rect 158078 105814 158130 105866
rect 158130 105814 158132 105866
rect 158076 105812 158132 105814
rect 158180 105866 158236 105868
rect 158180 105814 158182 105866
rect 158182 105814 158234 105866
rect 158234 105814 158236 105866
rect 158180 105812 158236 105814
rect 158284 105866 158340 105868
rect 158284 105814 158286 105866
rect 158286 105814 158338 105866
rect 158338 105814 158340 105866
rect 158284 105812 158340 105814
rect 173436 105082 173492 105084
rect 173436 105030 173438 105082
rect 173438 105030 173490 105082
rect 173490 105030 173492 105082
rect 173436 105028 173492 105030
rect 173540 105082 173596 105084
rect 173540 105030 173542 105082
rect 173542 105030 173594 105082
rect 173594 105030 173596 105082
rect 173540 105028 173596 105030
rect 173644 105082 173700 105084
rect 173644 105030 173646 105082
rect 173646 105030 173698 105082
rect 173698 105030 173700 105082
rect 173644 105028 173700 105030
rect 158076 104298 158132 104300
rect 158076 104246 158078 104298
rect 158078 104246 158130 104298
rect 158130 104246 158132 104298
rect 158076 104244 158132 104246
rect 158180 104298 158236 104300
rect 158180 104246 158182 104298
rect 158182 104246 158234 104298
rect 158234 104246 158236 104298
rect 158180 104244 158236 104246
rect 158284 104298 158340 104300
rect 158284 104246 158286 104298
rect 158286 104246 158338 104298
rect 158338 104246 158340 104298
rect 158284 104244 158340 104246
rect 173436 103514 173492 103516
rect 173436 103462 173438 103514
rect 173438 103462 173490 103514
rect 173490 103462 173492 103514
rect 173436 103460 173492 103462
rect 173540 103514 173596 103516
rect 173540 103462 173542 103514
rect 173542 103462 173594 103514
rect 173594 103462 173596 103514
rect 173540 103460 173596 103462
rect 173644 103514 173700 103516
rect 173644 103462 173646 103514
rect 173646 103462 173698 103514
rect 173698 103462 173700 103514
rect 173644 103460 173700 103462
rect 158076 102730 158132 102732
rect 158076 102678 158078 102730
rect 158078 102678 158130 102730
rect 158130 102678 158132 102730
rect 158076 102676 158132 102678
rect 158180 102730 158236 102732
rect 158180 102678 158182 102730
rect 158182 102678 158234 102730
rect 158234 102678 158236 102730
rect 158180 102676 158236 102678
rect 158284 102730 158340 102732
rect 158284 102678 158286 102730
rect 158286 102678 158338 102730
rect 158338 102678 158340 102730
rect 158284 102676 158340 102678
rect 173436 101946 173492 101948
rect 173436 101894 173438 101946
rect 173438 101894 173490 101946
rect 173490 101894 173492 101946
rect 173436 101892 173492 101894
rect 173540 101946 173596 101948
rect 173540 101894 173542 101946
rect 173542 101894 173594 101946
rect 173594 101894 173596 101946
rect 173540 101892 173596 101894
rect 173644 101946 173700 101948
rect 173644 101894 173646 101946
rect 173646 101894 173698 101946
rect 173698 101894 173700 101946
rect 173644 101892 173700 101894
rect 158076 101162 158132 101164
rect 158076 101110 158078 101162
rect 158078 101110 158130 101162
rect 158130 101110 158132 101162
rect 158076 101108 158132 101110
rect 158180 101162 158236 101164
rect 158180 101110 158182 101162
rect 158182 101110 158234 101162
rect 158234 101110 158236 101162
rect 158180 101108 158236 101110
rect 158284 101162 158340 101164
rect 158284 101110 158286 101162
rect 158286 101110 158338 101162
rect 158338 101110 158340 101162
rect 158284 101108 158340 101110
rect 173436 100378 173492 100380
rect 173436 100326 173438 100378
rect 173438 100326 173490 100378
rect 173490 100326 173492 100378
rect 173436 100324 173492 100326
rect 173540 100378 173596 100380
rect 173540 100326 173542 100378
rect 173542 100326 173594 100378
rect 173594 100326 173596 100378
rect 173540 100324 173596 100326
rect 173644 100378 173700 100380
rect 173644 100326 173646 100378
rect 173646 100326 173698 100378
rect 173698 100326 173700 100378
rect 173644 100324 173700 100326
rect 158076 99594 158132 99596
rect 158076 99542 158078 99594
rect 158078 99542 158130 99594
rect 158130 99542 158132 99594
rect 158076 99540 158132 99542
rect 158180 99594 158236 99596
rect 158180 99542 158182 99594
rect 158182 99542 158234 99594
rect 158234 99542 158236 99594
rect 158180 99540 158236 99542
rect 158284 99594 158340 99596
rect 158284 99542 158286 99594
rect 158286 99542 158338 99594
rect 158338 99542 158340 99594
rect 158284 99540 158340 99542
rect 173436 98810 173492 98812
rect 173436 98758 173438 98810
rect 173438 98758 173490 98810
rect 173490 98758 173492 98810
rect 173436 98756 173492 98758
rect 173540 98810 173596 98812
rect 173540 98758 173542 98810
rect 173542 98758 173594 98810
rect 173594 98758 173596 98810
rect 173540 98756 173596 98758
rect 173644 98810 173700 98812
rect 173644 98758 173646 98810
rect 173646 98758 173698 98810
rect 173698 98758 173700 98810
rect 173644 98756 173700 98758
rect 158076 98026 158132 98028
rect 158076 97974 158078 98026
rect 158078 97974 158130 98026
rect 158130 97974 158132 98026
rect 158076 97972 158132 97974
rect 158180 98026 158236 98028
rect 158180 97974 158182 98026
rect 158182 97974 158234 98026
rect 158234 97974 158236 98026
rect 158180 97972 158236 97974
rect 158284 98026 158340 98028
rect 158284 97974 158286 98026
rect 158286 97974 158338 98026
rect 158338 97974 158340 98026
rect 158284 97972 158340 97974
rect 173436 97242 173492 97244
rect 173436 97190 173438 97242
rect 173438 97190 173490 97242
rect 173490 97190 173492 97242
rect 173436 97188 173492 97190
rect 173540 97242 173596 97244
rect 173540 97190 173542 97242
rect 173542 97190 173594 97242
rect 173594 97190 173596 97242
rect 173540 97188 173596 97190
rect 173644 97242 173700 97244
rect 173644 97190 173646 97242
rect 173646 97190 173698 97242
rect 173698 97190 173700 97242
rect 173644 97188 173700 97190
rect 158076 96458 158132 96460
rect 158076 96406 158078 96458
rect 158078 96406 158130 96458
rect 158130 96406 158132 96458
rect 158076 96404 158132 96406
rect 158180 96458 158236 96460
rect 158180 96406 158182 96458
rect 158182 96406 158234 96458
rect 158234 96406 158236 96458
rect 158180 96404 158236 96406
rect 158284 96458 158340 96460
rect 158284 96406 158286 96458
rect 158286 96406 158338 96458
rect 158338 96406 158340 96458
rect 158284 96404 158340 96406
rect 173436 95674 173492 95676
rect 173436 95622 173438 95674
rect 173438 95622 173490 95674
rect 173490 95622 173492 95674
rect 173436 95620 173492 95622
rect 173540 95674 173596 95676
rect 173540 95622 173542 95674
rect 173542 95622 173594 95674
rect 173594 95622 173596 95674
rect 173540 95620 173596 95622
rect 173644 95674 173700 95676
rect 173644 95622 173646 95674
rect 173646 95622 173698 95674
rect 173698 95622 173700 95674
rect 173644 95620 173700 95622
rect 158076 94890 158132 94892
rect 158076 94838 158078 94890
rect 158078 94838 158130 94890
rect 158130 94838 158132 94890
rect 158076 94836 158132 94838
rect 158180 94890 158236 94892
rect 158180 94838 158182 94890
rect 158182 94838 158234 94890
rect 158234 94838 158236 94890
rect 158180 94836 158236 94838
rect 158284 94890 158340 94892
rect 158284 94838 158286 94890
rect 158286 94838 158338 94890
rect 158338 94838 158340 94890
rect 158284 94836 158340 94838
rect 173436 94106 173492 94108
rect 173436 94054 173438 94106
rect 173438 94054 173490 94106
rect 173490 94054 173492 94106
rect 173436 94052 173492 94054
rect 173540 94106 173596 94108
rect 173540 94054 173542 94106
rect 173542 94054 173594 94106
rect 173594 94054 173596 94106
rect 173540 94052 173596 94054
rect 173644 94106 173700 94108
rect 173644 94054 173646 94106
rect 173646 94054 173698 94106
rect 173698 94054 173700 94106
rect 173644 94052 173700 94054
rect 158076 93322 158132 93324
rect 158076 93270 158078 93322
rect 158078 93270 158130 93322
rect 158130 93270 158132 93322
rect 158076 93268 158132 93270
rect 158180 93322 158236 93324
rect 158180 93270 158182 93322
rect 158182 93270 158234 93322
rect 158234 93270 158236 93322
rect 158180 93268 158236 93270
rect 158284 93322 158340 93324
rect 158284 93270 158286 93322
rect 158286 93270 158338 93322
rect 158338 93270 158340 93322
rect 158284 93268 158340 93270
rect 173436 92538 173492 92540
rect 173436 92486 173438 92538
rect 173438 92486 173490 92538
rect 173490 92486 173492 92538
rect 173436 92484 173492 92486
rect 173540 92538 173596 92540
rect 173540 92486 173542 92538
rect 173542 92486 173594 92538
rect 173594 92486 173596 92538
rect 173540 92484 173596 92486
rect 173644 92538 173700 92540
rect 173644 92486 173646 92538
rect 173646 92486 173698 92538
rect 173698 92486 173700 92538
rect 173644 92484 173700 92486
rect 158076 91754 158132 91756
rect 158076 91702 158078 91754
rect 158078 91702 158130 91754
rect 158130 91702 158132 91754
rect 158076 91700 158132 91702
rect 158180 91754 158236 91756
rect 158180 91702 158182 91754
rect 158182 91702 158234 91754
rect 158234 91702 158236 91754
rect 158180 91700 158236 91702
rect 158284 91754 158340 91756
rect 158284 91702 158286 91754
rect 158286 91702 158338 91754
rect 158338 91702 158340 91754
rect 158284 91700 158340 91702
rect 173436 90970 173492 90972
rect 173436 90918 173438 90970
rect 173438 90918 173490 90970
rect 173490 90918 173492 90970
rect 173436 90916 173492 90918
rect 173540 90970 173596 90972
rect 173540 90918 173542 90970
rect 173542 90918 173594 90970
rect 173594 90918 173596 90970
rect 173540 90916 173596 90918
rect 173644 90970 173700 90972
rect 173644 90918 173646 90970
rect 173646 90918 173698 90970
rect 173698 90918 173700 90970
rect 173644 90916 173700 90918
rect 158076 90186 158132 90188
rect 158076 90134 158078 90186
rect 158078 90134 158130 90186
rect 158130 90134 158132 90186
rect 158076 90132 158132 90134
rect 158180 90186 158236 90188
rect 158180 90134 158182 90186
rect 158182 90134 158234 90186
rect 158234 90134 158236 90186
rect 158180 90132 158236 90134
rect 158284 90186 158340 90188
rect 158284 90134 158286 90186
rect 158286 90134 158338 90186
rect 158338 90134 158340 90186
rect 158284 90132 158340 90134
rect 173436 89402 173492 89404
rect 173436 89350 173438 89402
rect 173438 89350 173490 89402
rect 173490 89350 173492 89402
rect 173436 89348 173492 89350
rect 173540 89402 173596 89404
rect 173540 89350 173542 89402
rect 173542 89350 173594 89402
rect 173594 89350 173596 89402
rect 173540 89348 173596 89350
rect 173644 89402 173700 89404
rect 173644 89350 173646 89402
rect 173646 89350 173698 89402
rect 173698 89350 173700 89402
rect 173644 89348 173700 89350
rect 158076 88618 158132 88620
rect 158076 88566 158078 88618
rect 158078 88566 158130 88618
rect 158130 88566 158132 88618
rect 158076 88564 158132 88566
rect 158180 88618 158236 88620
rect 158180 88566 158182 88618
rect 158182 88566 158234 88618
rect 158234 88566 158236 88618
rect 158180 88564 158236 88566
rect 158284 88618 158340 88620
rect 158284 88566 158286 88618
rect 158286 88566 158338 88618
rect 158338 88566 158340 88618
rect 158284 88564 158340 88566
rect 173436 87834 173492 87836
rect 173436 87782 173438 87834
rect 173438 87782 173490 87834
rect 173490 87782 173492 87834
rect 173436 87780 173492 87782
rect 173540 87834 173596 87836
rect 173540 87782 173542 87834
rect 173542 87782 173594 87834
rect 173594 87782 173596 87834
rect 173540 87780 173596 87782
rect 173644 87834 173700 87836
rect 173644 87782 173646 87834
rect 173646 87782 173698 87834
rect 173698 87782 173700 87834
rect 173644 87780 173700 87782
rect 158076 87050 158132 87052
rect 158076 86998 158078 87050
rect 158078 86998 158130 87050
rect 158130 86998 158132 87050
rect 158076 86996 158132 86998
rect 158180 87050 158236 87052
rect 158180 86998 158182 87050
rect 158182 86998 158234 87050
rect 158234 86998 158236 87050
rect 158180 86996 158236 86998
rect 158284 87050 158340 87052
rect 158284 86998 158286 87050
rect 158286 86998 158338 87050
rect 158338 86998 158340 87050
rect 158284 86996 158340 86998
rect 173436 86266 173492 86268
rect 173436 86214 173438 86266
rect 173438 86214 173490 86266
rect 173490 86214 173492 86266
rect 173436 86212 173492 86214
rect 173540 86266 173596 86268
rect 173540 86214 173542 86266
rect 173542 86214 173594 86266
rect 173594 86214 173596 86266
rect 173540 86212 173596 86214
rect 173644 86266 173700 86268
rect 173644 86214 173646 86266
rect 173646 86214 173698 86266
rect 173698 86214 173700 86266
rect 173644 86212 173700 86214
rect 158076 85482 158132 85484
rect 158076 85430 158078 85482
rect 158078 85430 158130 85482
rect 158130 85430 158132 85482
rect 158076 85428 158132 85430
rect 158180 85482 158236 85484
rect 158180 85430 158182 85482
rect 158182 85430 158234 85482
rect 158234 85430 158236 85482
rect 158180 85428 158236 85430
rect 158284 85482 158340 85484
rect 158284 85430 158286 85482
rect 158286 85430 158338 85482
rect 158338 85430 158340 85482
rect 158284 85428 158340 85430
rect 173436 84698 173492 84700
rect 173436 84646 173438 84698
rect 173438 84646 173490 84698
rect 173490 84646 173492 84698
rect 173436 84644 173492 84646
rect 173540 84698 173596 84700
rect 173540 84646 173542 84698
rect 173542 84646 173594 84698
rect 173594 84646 173596 84698
rect 173540 84644 173596 84646
rect 173644 84698 173700 84700
rect 173644 84646 173646 84698
rect 173646 84646 173698 84698
rect 173698 84646 173700 84698
rect 173644 84644 173700 84646
rect 158076 83914 158132 83916
rect 158076 83862 158078 83914
rect 158078 83862 158130 83914
rect 158130 83862 158132 83914
rect 158076 83860 158132 83862
rect 158180 83914 158236 83916
rect 158180 83862 158182 83914
rect 158182 83862 158234 83914
rect 158234 83862 158236 83914
rect 158180 83860 158236 83862
rect 158284 83914 158340 83916
rect 158284 83862 158286 83914
rect 158286 83862 158338 83914
rect 158338 83862 158340 83914
rect 158284 83860 158340 83862
rect 173436 83130 173492 83132
rect 173436 83078 173438 83130
rect 173438 83078 173490 83130
rect 173490 83078 173492 83130
rect 173436 83076 173492 83078
rect 173540 83130 173596 83132
rect 173540 83078 173542 83130
rect 173542 83078 173594 83130
rect 173594 83078 173596 83130
rect 173540 83076 173596 83078
rect 173644 83130 173700 83132
rect 173644 83078 173646 83130
rect 173646 83078 173698 83130
rect 173698 83078 173700 83130
rect 173644 83076 173700 83078
rect 158076 82346 158132 82348
rect 158076 82294 158078 82346
rect 158078 82294 158130 82346
rect 158130 82294 158132 82346
rect 158076 82292 158132 82294
rect 158180 82346 158236 82348
rect 158180 82294 158182 82346
rect 158182 82294 158234 82346
rect 158234 82294 158236 82346
rect 158180 82292 158236 82294
rect 158284 82346 158340 82348
rect 158284 82294 158286 82346
rect 158286 82294 158338 82346
rect 158338 82294 158340 82346
rect 158284 82292 158340 82294
rect 173436 81562 173492 81564
rect 173436 81510 173438 81562
rect 173438 81510 173490 81562
rect 173490 81510 173492 81562
rect 173436 81508 173492 81510
rect 173540 81562 173596 81564
rect 173540 81510 173542 81562
rect 173542 81510 173594 81562
rect 173594 81510 173596 81562
rect 173540 81508 173596 81510
rect 173644 81562 173700 81564
rect 173644 81510 173646 81562
rect 173646 81510 173698 81562
rect 173698 81510 173700 81562
rect 173644 81508 173700 81510
rect 158076 80778 158132 80780
rect 158076 80726 158078 80778
rect 158078 80726 158130 80778
rect 158130 80726 158132 80778
rect 158076 80724 158132 80726
rect 158180 80778 158236 80780
rect 158180 80726 158182 80778
rect 158182 80726 158234 80778
rect 158234 80726 158236 80778
rect 158180 80724 158236 80726
rect 158284 80778 158340 80780
rect 158284 80726 158286 80778
rect 158286 80726 158338 80778
rect 158338 80726 158340 80778
rect 158284 80724 158340 80726
rect 173436 79994 173492 79996
rect 173436 79942 173438 79994
rect 173438 79942 173490 79994
rect 173490 79942 173492 79994
rect 173436 79940 173492 79942
rect 173540 79994 173596 79996
rect 173540 79942 173542 79994
rect 173542 79942 173594 79994
rect 173594 79942 173596 79994
rect 173540 79940 173596 79942
rect 173644 79994 173700 79996
rect 173644 79942 173646 79994
rect 173646 79942 173698 79994
rect 173698 79942 173700 79994
rect 173644 79940 173700 79942
rect 158076 79210 158132 79212
rect 158076 79158 158078 79210
rect 158078 79158 158130 79210
rect 158130 79158 158132 79210
rect 158076 79156 158132 79158
rect 158180 79210 158236 79212
rect 158180 79158 158182 79210
rect 158182 79158 158234 79210
rect 158234 79158 158236 79210
rect 158180 79156 158236 79158
rect 158284 79210 158340 79212
rect 158284 79158 158286 79210
rect 158286 79158 158338 79210
rect 158338 79158 158340 79210
rect 158284 79156 158340 79158
rect 173436 78426 173492 78428
rect 173436 78374 173438 78426
rect 173438 78374 173490 78426
rect 173490 78374 173492 78426
rect 173436 78372 173492 78374
rect 173540 78426 173596 78428
rect 173540 78374 173542 78426
rect 173542 78374 173594 78426
rect 173594 78374 173596 78426
rect 173540 78372 173596 78374
rect 173644 78426 173700 78428
rect 173644 78374 173646 78426
rect 173646 78374 173698 78426
rect 173698 78374 173700 78426
rect 173644 78372 173700 78374
rect 158076 77642 158132 77644
rect 158076 77590 158078 77642
rect 158078 77590 158130 77642
rect 158130 77590 158132 77642
rect 158076 77588 158132 77590
rect 158180 77642 158236 77644
rect 158180 77590 158182 77642
rect 158182 77590 158234 77642
rect 158234 77590 158236 77642
rect 158180 77588 158236 77590
rect 158284 77642 158340 77644
rect 158284 77590 158286 77642
rect 158286 77590 158338 77642
rect 158338 77590 158340 77642
rect 158284 77588 158340 77590
rect 173436 76858 173492 76860
rect 173436 76806 173438 76858
rect 173438 76806 173490 76858
rect 173490 76806 173492 76858
rect 173436 76804 173492 76806
rect 173540 76858 173596 76860
rect 173540 76806 173542 76858
rect 173542 76806 173594 76858
rect 173594 76806 173596 76858
rect 173540 76804 173596 76806
rect 173644 76858 173700 76860
rect 173644 76806 173646 76858
rect 173646 76806 173698 76858
rect 173698 76806 173700 76858
rect 173644 76804 173700 76806
rect 158076 76074 158132 76076
rect 158076 76022 158078 76074
rect 158078 76022 158130 76074
rect 158130 76022 158132 76074
rect 158076 76020 158132 76022
rect 158180 76074 158236 76076
rect 158180 76022 158182 76074
rect 158182 76022 158234 76074
rect 158234 76022 158236 76074
rect 158180 76020 158236 76022
rect 158284 76074 158340 76076
rect 158284 76022 158286 76074
rect 158286 76022 158338 76074
rect 158338 76022 158340 76074
rect 158284 76020 158340 76022
rect 173436 75290 173492 75292
rect 173436 75238 173438 75290
rect 173438 75238 173490 75290
rect 173490 75238 173492 75290
rect 173436 75236 173492 75238
rect 173540 75290 173596 75292
rect 173540 75238 173542 75290
rect 173542 75238 173594 75290
rect 173594 75238 173596 75290
rect 173540 75236 173596 75238
rect 173644 75290 173700 75292
rect 173644 75238 173646 75290
rect 173646 75238 173698 75290
rect 173698 75238 173700 75290
rect 173644 75236 173700 75238
rect 158076 74506 158132 74508
rect 158076 74454 158078 74506
rect 158078 74454 158130 74506
rect 158130 74454 158132 74506
rect 158076 74452 158132 74454
rect 158180 74506 158236 74508
rect 158180 74454 158182 74506
rect 158182 74454 158234 74506
rect 158234 74454 158236 74506
rect 158180 74452 158236 74454
rect 158284 74506 158340 74508
rect 158284 74454 158286 74506
rect 158286 74454 158338 74506
rect 158338 74454 158340 74506
rect 158284 74452 158340 74454
rect 173436 73722 173492 73724
rect 173436 73670 173438 73722
rect 173438 73670 173490 73722
rect 173490 73670 173492 73722
rect 173436 73668 173492 73670
rect 173540 73722 173596 73724
rect 173540 73670 173542 73722
rect 173542 73670 173594 73722
rect 173594 73670 173596 73722
rect 173540 73668 173596 73670
rect 173644 73722 173700 73724
rect 173644 73670 173646 73722
rect 173646 73670 173698 73722
rect 173698 73670 173700 73722
rect 173644 73668 173700 73670
rect 158076 72938 158132 72940
rect 158076 72886 158078 72938
rect 158078 72886 158130 72938
rect 158130 72886 158132 72938
rect 158076 72884 158132 72886
rect 158180 72938 158236 72940
rect 158180 72886 158182 72938
rect 158182 72886 158234 72938
rect 158234 72886 158236 72938
rect 158180 72884 158236 72886
rect 158284 72938 158340 72940
rect 158284 72886 158286 72938
rect 158286 72886 158338 72938
rect 158338 72886 158340 72938
rect 158284 72884 158340 72886
rect 173436 72154 173492 72156
rect 173436 72102 173438 72154
rect 173438 72102 173490 72154
rect 173490 72102 173492 72154
rect 173436 72100 173492 72102
rect 173540 72154 173596 72156
rect 173540 72102 173542 72154
rect 173542 72102 173594 72154
rect 173594 72102 173596 72154
rect 173540 72100 173596 72102
rect 173644 72154 173700 72156
rect 173644 72102 173646 72154
rect 173646 72102 173698 72154
rect 173698 72102 173700 72154
rect 173644 72100 173700 72102
rect 158076 71370 158132 71372
rect 158076 71318 158078 71370
rect 158078 71318 158130 71370
rect 158130 71318 158132 71370
rect 158076 71316 158132 71318
rect 158180 71370 158236 71372
rect 158180 71318 158182 71370
rect 158182 71318 158234 71370
rect 158234 71318 158236 71370
rect 158180 71316 158236 71318
rect 158284 71370 158340 71372
rect 158284 71318 158286 71370
rect 158286 71318 158338 71370
rect 158338 71318 158340 71370
rect 158284 71316 158340 71318
rect 173436 70586 173492 70588
rect 173436 70534 173438 70586
rect 173438 70534 173490 70586
rect 173490 70534 173492 70586
rect 173436 70532 173492 70534
rect 173540 70586 173596 70588
rect 173540 70534 173542 70586
rect 173542 70534 173594 70586
rect 173594 70534 173596 70586
rect 173540 70532 173596 70534
rect 173644 70586 173700 70588
rect 173644 70534 173646 70586
rect 173646 70534 173698 70586
rect 173698 70534 173700 70586
rect 173644 70532 173700 70534
rect 158076 69802 158132 69804
rect 158076 69750 158078 69802
rect 158078 69750 158130 69802
rect 158130 69750 158132 69802
rect 158076 69748 158132 69750
rect 158180 69802 158236 69804
rect 158180 69750 158182 69802
rect 158182 69750 158234 69802
rect 158234 69750 158236 69802
rect 158180 69748 158236 69750
rect 158284 69802 158340 69804
rect 158284 69750 158286 69802
rect 158286 69750 158338 69802
rect 158338 69750 158340 69802
rect 158284 69748 158340 69750
rect 173436 69018 173492 69020
rect 173436 68966 173438 69018
rect 173438 68966 173490 69018
rect 173490 68966 173492 69018
rect 173436 68964 173492 68966
rect 173540 69018 173596 69020
rect 173540 68966 173542 69018
rect 173542 68966 173594 69018
rect 173594 68966 173596 69018
rect 173540 68964 173596 68966
rect 173644 69018 173700 69020
rect 173644 68966 173646 69018
rect 173646 68966 173698 69018
rect 173698 68966 173700 69018
rect 173644 68964 173700 68966
rect 158076 68234 158132 68236
rect 158076 68182 158078 68234
rect 158078 68182 158130 68234
rect 158130 68182 158132 68234
rect 158076 68180 158132 68182
rect 158180 68234 158236 68236
rect 158180 68182 158182 68234
rect 158182 68182 158234 68234
rect 158234 68182 158236 68234
rect 158180 68180 158236 68182
rect 158284 68234 158340 68236
rect 158284 68182 158286 68234
rect 158286 68182 158338 68234
rect 158338 68182 158340 68234
rect 158284 68180 158340 68182
rect 173436 67450 173492 67452
rect 173436 67398 173438 67450
rect 173438 67398 173490 67450
rect 173490 67398 173492 67450
rect 173436 67396 173492 67398
rect 173540 67450 173596 67452
rect 173540 67398 173542 67450
rect 173542 67398 173594 67450
rect 173594 67398 173596 67450
rect 173540 67396 173596 67398
rect 173644 67450 173700 67452
rect 173644 67398 173646 67450
rect 173646 67398 173698 67450
rect 173698 67398 173700 67450
rect 173644 67396 173700 67398
rect 158076 66666 158132 66668
rect 158076 66614 158078 66666
rect 158078 66614 158130 66666
rect 158130 66614 158132 66666
rect 158076 66612 158132 66614
rect 158180 66666 158236 66668
rect 158180 66614 158182 66666
rect 158182 66614 158234 66666
rect 158234 66614 158236 66666
rect 158180 66612 158236 66614
rect 158284 66666 158340 66668
rect 158284 66614 158286 66666
rect 158286 66614 158338 66666
rect 158338 66614 158340 66666
rect 158284 66612 158340 66614
rect 173436 65882 173492 65884
rect 173436 65830 173438 65882
rect 173438 65830 173490 65882
rect 173490 65830 173492 65882
rect 173436 65828 173492 65830
rect 173540 65882 173596 65884
rect 173540 65830 173542 65882
rect 173542 65830 173594 65882
rect 173594 65830 173596 65882
rect 173540 65828 173596 65830
rect 173644 65882 173700 65884
rect 173644 65830 173646 65882
rect 173646 65830 173698 65882
rect 173698 65830 173700 65882
rect 173644 65828 173700 65830
rect 158076 65098 158132 65100
rect 158076 65046 158078 65098
rect 158078 65046 158130 65098
rect 158130 65046 158132 65098
rect 158076 65044 158132 65046
rect 158180 65098 158236 65100
rect 158180 65046 158182 65098
rect 158182 65046 158234 65098
rect 158234 65046 158236 65098
rect 158180 65044 158236 65046
rect 158284 65098 158340 65100
rect 158284 65046 158286 65098
rect 158286 65046 158338 65098
rect 158338 65046 158340 65098
rect 158284 65044 158340 65046
rect 173436 64314 173492 64316
rect 173436 64262 173438 64314
rect 173438 64262 173490 64314
rect 173490 64262 173492 64314
rect 173436 64260 173492 64262
rect 173540 64314 173596 64316
rect 173540 64262 173542 64314
rect 173542 64262 173594 64314
rect 173594 64262 173596 64314
rect 173540 64260 173596 64262
rect 173644 64314 173700 64316
rect 173644 64262 173646 64314
rect 173646 64262 173698 64314
rect 173698 64262 173700 64314
rect 173644 64260 173700 64262
rect 158076 63530 158132 63532
rect 158076 63478 158078 63530
rect 158078 63478 158130 63530
rect 158130 63478 158132 63530
rect 158076 63476 158132 63478
rect 158180 63530 158236 63532
rect 158180 63478 158182 63530
rect 158182 63478 158234 63530
rect 158234 63478 158236 63530
rect 158180 63476 158236 63478
rect 158284 63530 158340 63532
rect 158284 63478 158286 63530
rect 158286 63478 158338 63530
rect 158338 63478 158340 63530
rect 158284 63476 158340 63478
rect 173436 62746 173492 62748
rect 173436 62694 173438 62746
rect 173438 62694 173490 62746
rect 173490 62694 173492 62746
rect 173436 62692 173492 62694
rect 173540 62746 173596 62748
rect 173540 62694 173542 62746
rect 173542 62694 173594 62746
rect 173594 62694 173596 62746
rect 173540 62692 173596 62694
rect 173644 62746 173700 62748
rect 173644 62694 173646 62746
rect 173646 62694 173698 62746
rect 173698 62694 173700 62746
rect 173644 62692 173700 62694
rect 158076 61962 158132 61964
rect 158076 61910 158078 61962
rect 158078 61910 158130 61962
rect 158130 61910 158132 61962
rect 158076 61908 158132 61910
rect 158180 61962 158236 61964
rect 158180 61910 158182 61962
rect 158182 61910 158234 61962
rect 158234 61910 158236 61962
rect 158180 61908 158236 61910
rect 158284 61962 158340 61964
rect 158284 61910 158286 61962
rect 158286 61910 158338 61962
rect 158338 61910 158340 61962
rect 158284 61908 158340 61910
rect 173436 61178 173492 61180
rect 173436 61126 173438 61178
rect 173438 61126 173490 61178
rect 173490 61126 173492 61178
rect 173436 61124 173492 61126
rect 173540 61178 173596 61180
rect 173540 61126 173542 61178
rect 173542 61126 173594 61178
rect 173594 61126 173596 61178
rect 173540 61124 173596 61126
rect 173644 61178 173700 61180
rect 173644 61126 173646 61178
rect 173646 61126 173698 61178
rect 173698 61126 173700 61178
rect 173644 61124 173700 61126
rect 158076 60394 158132 60396
rect 158076 60342 158078 60394
rect 158078 60342 158130 60394
rect 158130 60342 158132 60394
rect 158076 60340 158132 60342
rect 158180 60394 158236 60396
rect 158180 60342 158182 60394
rect 158182 60342 158234 60394
rect 158234 60342 158236 60394
rect 158180 60340 158236 60342
rect 158284 60394 158340 60396
rect 158284 60342 158286 60394
rect 158286 60342 158338 60394
rect 158338 60342 158340 60394
rect 158284 60340 158340 60342
rect 173436 59610 173492 59612
rect 173436 59558 173438 59610
rect 173438 59558 173490 59610
rect 173490 59558 173492 59610
rect 173436 59556 173492 59558
rect 173540 59610 173596 59612
rect 173540 59558 173542 59610
rect 173542 59558 173594 59610
rect 173594 59558 173596 59610
rect 173540 59556 173596 59558
rect 173644 59610 173700 59612
rect 173644 59558 173646 59610
rect 173646 59558 173698 59610
rect 173698 59558 173700 59610
rect 173644 59556 173700 59558
rect 158076 58826 158132 58828
rect 158076 58774 158078 58826
rect 158078 58774 158130 58826
rect 158130 58774 158132 58826
rect 158076 58772 158132 58774
rect 158180 58826 158236 58828
rect 158180 58774 158182 58826
rect 158182 58774 158234 58826
rect 158234 58774 158236 58826
rect 158180 58772 158236 58774
rect 158284 58826 158340 58828
rect 158284 58774 158286 58826
rect 158286 58774 158338 58826
rect 158338 58774 158340 58826
rect 158284 58772 158340 58774
rect 173436 58042 173492 58044
rect 173436 57990 173438 58042
rect 173438 57990 173490 58042
rect 173490 57990 173492 58042
rect 173436 57988 173492 57990
rect 173540 58042 173596 58044
rect 173540 57990 173542 58042
rect 173542 57990 173594 58042
rect 173594 57990 173596 58042
rect 173540 57988 173596 57990
rect 173644 58042 173700 58044
rect 173644 57990 173646 58042
rect 173646 57990 173698 58042
rect 173698 57990 173700 58042
rect 173644 57988 173700 57990
rect 158076 57258 158132 57260
rect 158076 57206 158078 57258
rect 158078 57206 158130 57258
rect 158130 57206 158132 57258
rect 158076 57204 158132 57206
rect 158180 57258 158236 57260
rect 158180 57206 158182 57258
rect 158182 57206 158234 57258
rect 158234 57206 158236 57258
rect 158180 57204 158236 57206
rect 158284 57258 158340 57260
rect 158284 57206 158286 57258
rect 158286 57206 158338 57258
rect 158338 57206 158340 57258
rect 158284 57204 158340 57206
rect 173436 56474 173492 56476
rect 173436 56422 173438 56474
rect 173438 56422 173490 56474
rect 173490 56422 173492 56474
rect 173436 56420 173492 56422
rect 173540 56474 173596 56476
rect 173540 56422 173542 56474
rect 173542 56422 173594 56474
rect 173594 56422 173596 56474
rect 173540 56420 173596 56422
rect 173644 56474 173700 56476
rect 173644 56422 173646 56474
rect 173646 56422 173698 56474
rect 173698 56422 173700 56474
rect 173644 56420 173700 56422
rect 158076 55690 158132 55692
rect 158076 55638 158078 55690
rect 158078 55638 158130 55690
rect 158130 55638 158132 55690
rect 158076 55636 158132 55638
rect 158180 55690 158236 55692
rect 158180 55638 158182 55690
rect 158182 55638 158234 55690
rect 158234 55638 158236 55690
rect 158180 55636 158236 55638
rect 158284 55690 158340 55692
rect 158284 55638 158286 55690
rect 158286 55638 158338 55690
rect 158338 55638 158340 55690
rect 158284 55636 158340 55638
rect 173436 54906 173492 54908
rect 173436 54854 173438 54906
rect 173438 54854 173490 54906
rect 173490 54854 173492 54906
rect 173436 54852 173492 54854
rect 173540 54906 173596 54908
rect 173540 54854 173542 54906
rect 173542 54854 173594 54906
rect 173594 54854 173596 54906
rect 173540 54852 173596 54854
rect 173644 54906 173700 54908
rect 173644 54854 173646 54906
rect 173646 54854 173698 54906
rect 173698 54854 173700 54906
rect 173644 54852 173700 54854
rect 158076 54122 158132 54124
rect 158076 54070 158078 54122
rect 158078 54070 158130 54122
rect 158130 54070 158132 54122
rect 158076 54068 158132 54070
rect 158180 54122 158236 54124
rect 158180 54070 158182 54122
rect 158182 54070 158234 54122
rect 158234 54070 158236 54122
rect 158180 54068 158236 54070
rect 158284 54122 158340 54124
rect 158284 54070 158286 54122
rect 158286 54070 158338 54122
rect 158338 54070 158340 54122
rect 158284 54068 158340 54070
rect 173436 53338 173492 53340
rect 173436 53286 173438 53338
rect 173438 53286 173490 53338
rect 173490 53286 173492 53338
rect 173436 53284 173492 53286
rect 173540 53338 173596 53340
rect 173540 53286 173542 53338
rect 173542 53286 173594 53338
rect 173594 53286 173596 53338
rect 173540 53284 173596 53286
rect 173644 53338 173700 53340
rect 173644 53286 173646 53338
rect 173646 53286 173698 53338
rect 173698 53286 173700 53338
rect 173644 53284 173700 53286
rect 158076 52554 158132 52556
rect 158076 52502 158078 52554
rect 158078 52502 158130 52554
rect 158130 52502 158132 52554
rect 158076 52500 158132 52502
rect 158180 52554 158236 52556
rect 158180 52502 158182 52554
rect 158182 52502 158234 52554
rect 158234 52502 158236 52554
rect 158180 52500 158236 52502
rect 158284 52554 158340 52556
rect 158284 52502 158286 52554
rect 158286 52502 158338 52554
rect 158338 52502 158340 52554
rect 158284 52500 158340 52502
rect 173436 51770 173492 51772
rect 173436 51718 173438 51770
rect 173438 51718 173490 51770
rect 173490 51718 173492 51770
rect 173436 51716 173492 51718
rect 173540 51770 173596 51772
rect 173540 51718 173542 51770
rect 173542 51718 173594 51770
rect 173594 51718 173596 51770
rect 173540 51716 173596 51718
rect 173644 51770 173700 51772
rect 173644 51718 173646 51770
rect 173646 51718 173698 51770
rect 173698 51718 173700 51770
rect 173644 51716 173700 51718
rect 158076 50986 158132 50988
rect 158076 50934 158078 50986
rect 158078 50934 158130 50986
rect 158130 50934 158132 50986
rect 158076 50932 158132 50934
rect 158180 50986 158236 50988
rect 158180 50934 158182 50986
rect 158182 50934 158234 50986
rect 158234 50934 158236 50986
rect 158180 50932 158236 50934
rect 158284 50986 158340 50988
rect 158284 50934 158286 50986
rect 158286 50934 158338 50986
rect 158338 50934 158340 50986
rect 158284 50932 158340 50934
rect 173436 50202 173492 50204
rect 173436 50150 173438 50202
rect 173438 50150 173490 50202
rect 173490 50150 173492 50202
rect 173436 50148 173492 50150
rect 173540 50202 173596 50204
rect 173540 50150 173542 50202
rect 173542 50150 173594 50202
rect 173594 50150 173596 50202
rect 173540 50148 173596 50150
rect 173644 50202 173700 50204
rect 173644 50150 173646 50202
rect 173646 50150 173698 50202
rect 173698 50150 173700 50202
rect 173644 50148 173700 50150
rect 158076 49418 158132 49420
rect 158076 49366 158078 49418
rect 158078 49366 158130 49418
rect 158130 49366 158132 49418
rect 158076 49364 158132 49366
rect 158180 49418 158236 49420
rect 158180 49366 158182 49418
rect 158182 49366 158234 49418
rect 158234 49366 158236 49418
rect 158180 49364 158236 49366
rect 158284 49418 158340 49420
rect 158284 49366 158286 49418
rect 158286 49366 158338 49418
rect 158338 49366 158340 49418
rect 158284 49364 158340 49366
rect 173436 48634 173492 48636
rect 173436 48582 173438 48634
rect 173438 48582 173490 48634
rect 173490 48582 173492 48634
rect 173436 48580 173492 48582
rect 173540 48634 173596 48636
rect 173540 48582 173542 48634
rect 173542 48582 173594 48634
rect 173594 48582 173596 48634
rect 173540 48580 173596 48582
rect 173644 48634 173700 48636
rect 173644 48582 173646 48634
rect 173646 48582 173698 48634
rect 173698 48582 173700 48634
rect 173644 48580 173700 48582
rect 158076 47850 158132 47852
rect 158076 47798 158078 47850
rect 158078 47798 158130 47850
rect 158130 47798 158132 47850
rect 158076 47796 158132 47798
rect 158180 47850 158236 47852
rect 158180 47798 158182 47850
rect 158182 47798 158234 47850
rect 158234 47798 158236 47850
rect 158180 47796 158236 47798
rect 158284 47850 158340 47852
rect 158284 47798 158286 47850
rect 158286 47798 158338 47850
rect 158338 47798 158340 47850
rect 158284 47796 158340 47798
rect 173436 47066 173492 47068
rect 173436 47014 173438 47066
rect 173438 47014 173490 47066
rect 173490 47014 173492 47066
rect 173436 47012 173492 47014
rect 173540 47066 173596 47068
rect 173540 47014 173542 47066
rect 173542 47014 173594 47066
rect 173594 47014 173596 47066
rect 173540 47012 173596 47014
rect 173644 47066 173700 47068
rect 173644 47014 173646 47066
rect 173646 47014 173698 47066
rect 173698 47014 173700 47066
rect 173644 47012 173700 47014
rect 158076 46282 158132 46284
rect 158076 46230 158078 46282
rect 158078 46230 158130 46282
rect 158130 46230 158132 46282
rect 158076 46228 158132 46230
rect 158180 46282 158236 46284
rect 158180 46230 158182 46282
rect 158182 46230 158234 46282
rect 158234 46230 158236 46282
rect 158180 46228 158236 46230
rect 158284 46282 158340 46284
rect 158284 46230 158286 46282
rect 158286 46230 158338 46282
rect 158338 46230 158340 46282
rect 158284 46228 158340 46230
rect 173436 45498 173492 45500
rect 173436 45446 173438 45498
rect 173438 45446 173490 45498
rect 173490 45446 173492 45498
rect 173436 45444 173492 45446
rect 173540 45498 173596 45500
rect 173540 45446 173542 45498
rect 173542 45446 173594 45498
rect 173594 45446 173596 45498
rect 173540 45444 173596 45446
rect 173644 45498 173700 45500
rect 173644 45446 173646 45498
rect 173646 45446 173698 45498
rect 173698 45446 173700 45498
rect 173644 45444 173700 45446
rect 158076 44714 158132 44716
rect 158076 44662 158078 44714
rect 158078 44662 158130 44714
rect 158130 44662 158132 44714
rect 158076 44660 158132 44662
rect 158180 44714 158236 44716
rect 158180 44662 158182 44714
rect 158182 44662 158234 44714
rect 158234 44662 158236 44714
rect 158180 44660 158236 44662
rect 158284 44714 158340 44716
rect 158284 44662 158286 44714
rect 158286 44662 158338 44714
rect 158338 44662 158340 44714
rect 158284 44660 158340 44662
rect 173436 43930 173492 43932
rect 173436 43878 173438 43930
rect 173438 43878 173490 43930
rect 173490 43878 173492 43930
rect 173436 43876 173492 43878
rect 173540 43930 173596 43932
rect 173540 43878 173542 43930
rect 173542 43878 173594 43930
rect 173594 43878 173596 43930
rect 173540 43876 173596 43878
rect 173644 43930 173700 43932
rect 173644 43878 173646 43930
rect 173646 43878 173698 43930
rect 173698 43878 173700 43930
rect 173644 43876 173700 43878
rect 158076 43146 158132 43148
rect 158076 43094 158078 43146
rect 158078 43094 158130 43146
rect 158130 43094 158132 43146
rect 158076 43092 158132 43094
rect 158180 43146 158236 43148
rect 158180 43094 158182 43146
rect 158182 43094 158234 43146
rect 158234 43094 158236 43146
rect 158180 43092 158236 43094
rect 158284 43146 158340 43148
rect 158284 43094 158286 43146
rect 158286 43094 158338 43146
rect 158338 43094 158340 43146
rect 158284 43092 158340 43094
rect 173436 42362 173492 42364
rect 173436 42310 173438 42362
rect 173438 42310 173490 42362
rect 173490 42310 173492 42362
rect 173436 42308 173492 42310
rect 173540 42362 173596 42364
rect 173540 42310 173542 42362
rect 173542 42310 173594 42362
rect 173594 42310 173596 42362
rect 173540 42308 173596 42310
rect 173644 42362 173700 42364
rect 173644 42310 173646 42362
rect 173646 42310 173698 42362
rect 173698 42310 173700 42362
rect 173644 42308 173700 42310
rect 158076 41578 158132 41580
rect 158076 41526 158078 41578
rect 158078 41526 158130 41578
rect 158130 41526 158132 41578
rect 158076 41524 158132 41526
rect 158180 41578 158236 41580
rect 158180 41526 158182 41578
rect 158182 41526 158234 41578
rect 158234 41526 158236 41578
rect 158180 41524 158236 41526
rect 158284 41578 158340 41580
rect 158284 41526 158286 41578
rect 158286 41526 158338 41578
rect 158338 41526 158340 41578
rect 158284 41524 158340 41526
rect 173436 40794 173492 40796
rect 173436 40742 173438 40794
rect 173438 40742 173490 40794
rect 173490 40742 173492 40794
rect 173436 40740 173492 40742
rect 173540 40794 173596 40796
rect 173540 40742 173542 40794
rect 173542 40742 173594 40794
rect 173594 40742 173596 40794
rect 173540 40740 173596 40742
rect 173644 40794 173700 40796
rect 173644 40742 173646 40794
rect 173646 40742 173698 40794
rect 173698 40742 173700 40794
rect 173644 40740 173700 40742
rect 158076 40010 158132 40012
rect 158076 39958 158078 40010
rect 158078 39958 158130 40010
rect 158130 39958 158132 40010
rect 158076 39956 158132 39958
rect 158180 40010 158236 40012
rect 158180 39958 158182 40010
rect 158182 39958 158234 40010
rect 158234 39958 158236 40010
rect 158180 39956 158236 39958
rect 158284 40010 158340 40012
rect 158284 39958 158286 40010
rect 158286 39958 158338 40010
rect 158338 39958 158340 40010
rect 158284 39956 158340 39958
rect 173436 39226 173492 39228
rect 173436 39174 173438 39226
rect 173438 39174 173490 39226
rect 173490 39174 173492 39226
rect 173436 39172 173492 39174
rect 173540 39226 173596 39228
rect 173540 39174 173542 39226
rect 173542 39174 173594 39226
rect 173594 39174 173596 39226
rect 173540 39172 173596 39174
rect 173644 39226 173700 39228
rect 173644 39174 173646 39226
rect 173646 39174 173698 39226
rect 173698 39174 173700 39226
rect 173644 39172 173700 39174
rect 158076 38442 158132 38444
rect 158076 38390 158078 38442
rect 158078 38390 158130 38442
rect 158130 38390 158132 38442
rect 158076 38388 158132 38390
rect 158180 38442 158236 38444
rect 158180 38390 158182 38442
rect 158182 38390 158234 38442
rect 158234 38390 158236 38442
rect 158180 38388 158236 38390
rect 158284 38442 158340 38444
rect 158284 38390 158286 38442
rect 158286 38390 158338 38442
rect 158338 38390 158340 38442
rect 158284 38388 158340 38390
rect 173436 37658 173492 37660
rect 173436 37606 173438 37658
rect 173438 37606 173490 37658
rect 173490 37606 173492 37658
rect 173436 37604 173492 37606
rect 173540 37658 173596 37660
rect 173540 37606 173542 37658
rect 173542 37606 173594 37658
rect 173594 37606 173596 37658
rect 173540 37604 173596 37606
rect 173644 37658 173700 37660
rect 173644 37606 173646 37658
rect 173646 37606 173698 37658
rect 173698 37606 173700 37658
rect 173644 37604 173700 37606
rect 158076 36874 158132 36876
rect 158076 36822 158078 36874
rect 158078 36822 158130 36874
rect 158130 36822 158132 36874
rect 158076 36820 158132 36822
rect 158180 36874 158236 36876
rect 158180 36822 158182 36874
rect 158182 36822 158234 36874
rect 158234 36822 158236 36874
rect 158180 36820 158236 36822
rect 158284 36874 158340 36876
rect 158284 36822 158286 36874
rect 158286 36822 158338 36874
rect 158338 36822 158340 36874
rect 158284 36820 158340 36822
rect 173436 36090 173492 36092
rect 173436 36038 173438 36090
rect 173438 36038 173490 36090
rect 173490 36038 173492 36090
rect 173436 36036 173492 36038
rect 173540 36090 173596 36092
rect 173540 36038 173542 36090
rect 173542 36038 173594 36090
rect 173594 36038 173596 36090
rect 173540 36036 173596 36038
rect 173644 36090 173700 36092
rect 173644 36038 173646 36090
rect 173646 36038 173698 36090
rect 173698 36038 173700 36090
rect 173644 36036 173700 36038
rect 158076 35306 158132 35308
rect 158076 35254 158078 35306
rect 158078 35254 158130 35306
rect 158130 35254 158132 35306
rect 158076 35252 158132 35254
rect 158180 35306 158236 35308
rect 158180 35254 158182 35306
rect 158182 35254 158234 35306
rect 158234 35254 158236 35306
rect 158180 35252 158236 35254
rect 158284 35306 158340 35308
rect 158284 35254 158286 35306
rect 158286 35254 158338 35306
rect 158338 35254 158340 35306
rect 158284 35252 158340 35254
rect 173436 34522 173492 34524
rect 173436 34470 173438 34522
rect 173438 34470 173490 34522
rect 173490 34470 173492 34522
rect 173436 34468 173492 34470
rect 173540 34522 173596 34524
rect 173540 34470 173542 34522
rect 173542 34470 173594 34522
rect 173594 34470 173596 34522
rect 173540 34468 173596 34470
rect 173644 34522 173700 34524
rect 173644 34470 173646 34522
rect 173646 34470 173698 34522
rect 173698 34470 173700 34522
rect 173644 34468 173700 34470
rect 158076 33738 158132 33740
rect 158076 33686 158078 33738
rect 158078 33686 158130 33738
rect 158130 33686 158132 33738
rect 158076 33684 158132 33686
rect 158180 33738 158236 33740
rect 158180 33686 158182 33738
rect 158182 33686 158234 33738
rect 158234 33686 158236 33738
rect 158180 33684 158236 33686
rect 158284 33738 158340 33740
rect 158284 33686 158286 33738
rect 158286 33686 158338 33738
rect 158338 33686 158340 33738
rect 158284 33684 158340 33686
rect 173436 32954 173492 32956
rect 173436 32902 173438 32954
rect 173438 32902 173490 32954
rect 173490 32902 173492 32954
rect 173436 32900 173492 32902
rect 173540 32954 173596 32956
rect 173540 32902 173542 32954
rect 173542 32902 173594 32954
rect 173594 32902 173596 32954
rect 173540 32900 173596 32902
rect 173644 32954 173700 32956
rect 173644 32902 173646 32954
rect 173646 32902 173698 32954
rect 173698 32902 173700 32954
rect 173644 32900 173700 32902
rect 158076 32170 158132 32172
rect 158076 32118 158078 32170
rect 158078 32118 158130 32170
rect 158130 32118 158132 32170
rect 158076 32116 158132 32118
rect 158180 32170 158236 32172
rect 158180 32118 158182 32170
rect 158182 32118 158234 32170
rect 158234 32118 158236 32170
rect 158180 32116 158236 32118
rect 158284 32170 158340 32172
rect 158284 32118 158286 32170
rect 158286 32118 158338 32170
rect 158338 32118 158340 32170
rect 158284 32116 158340 32118
rect 173436 31386 173492 31388
rect 173436 31334 173438 31386
rect 173438 31334 173490 31386
rect 173490 31334 173492 31386
rect 173436 31332 173492 31334
rect 173540 31386 173596 31388
rect 173540 31334 173542 31386
rect 173542 31334 173594 31386
rect 173594 31334 173596 31386
rect 173540 31332 173596 31334
rect 173644 31386 173700 31388
rect 173644 31334 173646 31386
rect 173646 31334 173698 31386
rect 173698 31334 173700 31386
rect 173644 31332 173700 31334
rect 158076 30602 158132 30604
rect 158076 30550 158078 30602
rect 158078 30550 158130 30602
rect 158130 30550 158132 30602
rect 158076 30548 158132 30550
rect 158180 30602 158236 30604
rect 158180 30550 158182 30602
rect 158182 30550 158234 30602
rect 158234 30550 158236 30602
rect 158180 30548 158236 30550
rect 158284 30602 158340 30604
rect 158284 30550 158286 30602
rect 158286 30550 158338 30602
rect 158338 30550 158340 30602
rect 158284 30548 158340 30550
rect 173436 29818 173492 29820
rect 173436 29766 173438 29818
rect 173438 29766 173490 29818
rect 173490 29766 173492 29818
rect 173436 29764 173492 29766
rect 173540 29818 173596 29820
rect 173540 29766 173542 29818
rect 173542 29766 173594 29818
rect 173594 29766 173596 29818
rect 173540 29764 173596 29766
rect 173644 29818 173700 29820
rect 173644 29766 173646 29818
rect 173646 29766 173698 29818
rect 173698 29766 173700 29818
rect 173644 29764 173700 29766
rect 158076 29034 158132 29036
rect 158076 28982 158078 29034
rect 158078 28982 158130 29034
rect 158130 28982 158132 29034
rect 158076 28980 158132 28982
rect 158180 29034 158236 29036
rect 158180 28982 158182 29034
rect 158182 28982 158234 29034
rect 158234 28982 158236 29034
rect 158180 28980 158236 28982
rect 158284 29034 158340 29036
rect 158284 28982 158286 29034
rect 158286 28982 158338 29034
rect 158338 28982 158340 29034
rect 158284 28980 158340 28982
rect 173436 28250 173492 28252
rect 173436 28198 173438 28250
rect 173438 28198 173490 28250
rect 173490 28198 173492 28250
rect 173436 28196 173492 28198
rect 173540 28250 173596 28252
rect 173540 28198 173542 28250
rect 173542 28198 173594 28250
rect 173594 28198 173596 28250
rect 173540 28196 173596 28198
rect 173644 28250 173700 28252
rect 173644 28198 173646 28250
rect 173646 28198 173698 28250
rect 173698 28198 173700 28250
rect 173644 28196 173700 28198
rect 158076 27466 158132 27468
rect 158076 27414 158078 27466
rect 158078 27414 158130 27466
rect 158130 27414 158132 27466
rect 158076 27412 158132 27414
rect 158180 27466 158236 27468
rect 158180 27414 158182 27466
rect 158182 27414 158234 27466
rect 158234 27414 158236 27466
rect 158180 27412 158236 27414
rect 158284 27466 158340 27468
rect 158284 27414 158286 27466
rect 158286 27414 158338 27466
rect 158338 27414 158340 27466
rect 158284 27412 158340 27414
rect 173436 26682 173492 26684
rect 173436 26630 173438 26682
rect 173438 26630 173490 26682
rect 173490 26630 173492 26682
rect 173436 26628 173492 26630
rect 173540 26682 173596 26684
rect 173540 26630 173542 26682
rect 173542 26630 173594 26682
rect 173594 26630 173596 26682
rect 173540 26628 173596 26630
rect 173644 26682 173700 26684
rect 173644 26630 173646 26682
rect 173646 26630 173698 26682
rect 173698 26630 173700 26682
rect 173644 26628 173700 26630
rect 158076 25898 158132 25900
rect 158076 25846 158078 25898
rect 158078 25846 158130 25898
rect 158130 25846 158132 25898
rect 158076 25844 158132 25846
rect 158180 25898 158236 25900
rect 158180 25846 158182 25898
rect 158182 25846 158234 25898
rect 158234 25846 158236 25898
rect 158180 25844 158236 25846
rect 158284 25898 158340 25900
rect 158284 25846 158286 25898
rect 158286 25846 158338 25898
rect 158338 25846 158340 25898
rect 158284 25844 158340 25846
rect 173436 25114 173492 25116
rect 173436 25062 173438 25114
rect 173438 25062 173490 25114
rect 173490 25062 173492 25114
rect 173436 25060 173492 25062
rect 173540 25114 173596 25116
rect 173540 25062 173542 25114
rect 173542 25062 173594 25114
rect 173594 25062 173596 25114
rect 173540 25060 173596 25062
rect 173644 25114 173700 25116
rect 173644 25062 173646 25114
rect 173646 25062 173698 25114
rect 173698 25062 173700 25114
rect 173644 25060 173700 25062
rect 169148 24444 169204 24500
rect 158076 24330 158132 24332
rect 158076 24278 158078 24330
rect 158078 24278 158130 24330
rect 158130 24278 158132 24330
rect 158076 24276 158132 24278
rect 158180 24330 158236 24332
rect 158180 24278 158182 24330
rect 158182 24278 158234 24330
rect 158234 24278 158236 24330
rect 158180 24276 158236 24278
rect 158284 24330 158340 24332
rect 158284 24278 158286 24330
rect 158286 24278 158338 24330
rect 158338 24278 158340 24330
rect 158284 24276 158340 24278
rect 158076 22762 158132 22764
rect 158076 22710 158078 22762
rect 158078 22710 158130 22762
rect 158130 22710 158132 22762
rect 158076 22708 158132 22710
rect 158180 22762 158236 22764
rect 158180 22710 158182 22762
rect 158182 22710 158234 22762
rect 158234 22710 158236 22762
rect 158180 22708 158236 22710
rect 158284 22762 158340 22764
rect 158284 22710 158286 22762
rect 158286 22710 158338 22762
rect 158338 22710 158340 22762
rect 158284 22708 158340 22710
rect 158076 21194 158132 21196
rect 158076 21142 158078 21194
rect 158078 21142 158130 21194
rect 158130 21142 158132 21194
rect 158076 21140 158132 21142
rect 158180 21194 158236 21196
rect 158180 21142 158182 21194
rect 158182 21142 158234 21194
rect 158234 21142 158236 21194
rect 158180 21140 158236 21142
rect 158284 21194 158340 21196
rect 158284 21142 158286 21194
rect 158286 21142 158338 21194
rect 158338 21142 158340 21194
rect 158284 21140 158340 21142
rect 167356 20860 167412 20916
rect 158076 19626 158132 19628
rect 158076 19574 158078 19626
rect 158078 19574 158130 19626
rect 158130 19574 158132 19626
rect 158076 19572 158132 19574
rect 158180 19626 158236 19628
rect 158180 19574 158182 19626
rect 158182 19574 158234 19626
rect 158234 19574 158236 19626
rect 158180 19572 158236 19574
rect 158284 19626 158340 19628
rect 158284 19574 158286 19626
rect 158286 19574 158338 19626
rect 158338 19574 158340 19626
rect 158284 19572 158340 19574
rect 163436 18508 163492 18564
rect 158076 18058 158132 18060
rect 158076 18006 158078 18058
rect 158078 18006 158130 18058
rect 158130 18006 158132 18058
rect 158076 18004 158132 18006
rect 158180 18058 158236 18060
rect 158180 18006 158182 18058
rect 158182 18006 158234 18058
rect 158234 18006 158236 18058
rect 158180 18004 158236 18006
rect 158284 18058 158340 18060
rect 158284 18006 158286 18058
rect 158286 18006 158338 18058
rect 158338 18006 158340 18058
rect 158284 18004 158340 18006
rect 158076 16490 158132 16492
rect 158076 16438 158078 16490
rect 158078 16438 158130 16490
rect 158130 16438 158132 16490
rect 158076 16436 158132 16438
rect 158180 16490 158236 16492
rect 158180 16438 158182 16490
rect 158182 16438 158234 16490
rect 158234 16438 158236 16490
rect 158180 16436 158236 16438
rect 158284 16490 158340 16492
rect 158284 16438 158286 16490
rect 158286 16438 158338 16490
rect 158338 16438 158340 16490
rect 158284 16436 158340 16438
rect 158076 14922 158132 14924
rect 158076 14870 158078 14922
rect 158078 14870 158130 14922
rect 158130 14870 158132 14922
rect 158076 14868 158132 14870
rect 158180 14922 158236 14924
rect 158180 14870 158182 14922
rect 158182 14870 158234 14922
rect 158234 14870 158236 14922
rect 158180 14868 158236 14870
rect 158284 14922 158340 14924
rect 158284 14870 158286 14922
rect 158286 14870 158338 14922
rect 158338 14870 158340 14922
rect 158284 14868 158340 14870
rect 161308 13580 161364 13636
rect 158076 13354 158132 13356
rect 158076 13302 158078 13354
rect 158078 13302 158130 13354
rect 158130 13302 158132 13354
rect 158076 13300 158132 13302
rect 158180 13354 158236 13356
rect 158180 13302 158182 13354
rect 158182 13302 158234 13354
rect 158234 13302 158236 13354
rect 158180 13300 158236 13302
rect 158284 13354 158340 13356
rect 158284 13302 158286 13354
rect 158286 13302 158338 13354
rect 158338 13302 158340 13354
rect 158284 13300 158340 13302
rect 158076 11786 158132 11788
rect 158076 11734 158078 11786
rect 158078 11734 158130 11786
rect 158130 11734 158132 11786
rect 158076 11732 158132 11734
rect 158180 11786 158236 11788
rect 158180 11734 158182 11786
rect 158182 11734 158234 11786
rect 158234 11734 158236 11786
rect 158180 11732 158236 11734
rect 158284 11786 158340 11788
rect 158284 11734 158286 11786
rect 158286 11734 158338 11786
rect 158338 11734 158340 11786
rect 158284 11732 158340 11734
rect 150444 11116 150500 11172
rect 160412 10780 160468 10836
rect 156268 10444 156324 10500
rect 148876 8988 148932 9044
rect 146076 5628 146132 5684
rect 146188 5010 146244 5012
rect 146188 4958 146190 5010
rect 146190 4958 146242 5010
rect 146242 4958 146244 5010
rect 146188 4956 146244 4958
rect 146636 6466 146692 6468
rect 146636 6414 146638 6466
rect 146638 6414 146690 6466
rect 146690 6414 146692 6466
rect 146636 6412 146692 6414
rect 146972 6412 147028 6468
rect 146300 3948 146356 4004
rect 145628 3724 145684 3780
rect 145292 3388 145348 3444
rect 145404 3500 145460 3556
rect 146076 3612 146132 3668
rect 145964 3442 146020 3444
rect 145964 3390 145966 3442
rect 145966 3390 146018 3442
rect 146018 3390 146020 3442
rect 145964 3388 146020 3390
rect 146748 5010 146804 5012
rect 146748 4958 146750 5010
rect 146750 4958 146802 5010
rect 146802 4958 146804 5010
rect 146748 4956 146804 4958
rect 147084 5180 147140 5236
rect 147308 5794 147364 5796
rect 147308 5742 147310 5794
rect 147310 5742 147362 5794
rect 147362 5742 147364 5794
rect 147308 5740 147364 5742
rect 147308 5292 147364 5348
rect 147308 4338 147364 4340
rect 147308 4286 147310 4338
rect 147310 4286 147362 4338
rect 147362 4286 147364 4338
rect 147308 4284 147364 4286
rect 147196 3554 147252 3556
rect 147196 3502 147198 3554
rect 147198 3502 147250 3554
rect 147250 3502 147252 3554
rect 147196 3500 147252 3502
rect 147084 3388 147140 3444
rect 146860 3330 146916 3332
rect 146860 3278 146862 3330
rect 146862 3278 146914 3330
rect 146914 3278 146916 3330
rect 146860 3276 146916 3278
rect 147644 5234 147700 5236
rect 147644 5182 147646 5234
rect 147646 5182 147698 5234
rect 147698 5182 147700 5234
rect 147644 5180 147700 5182
rect 147756 5010 147812 5012
rect 147756 4958 147758 5010
rect 147758 4958 147810 5010
rect 147810 4958 147812 5010
rect 147756 4956 147812 4958
rect 147532 3612 147588 3668
rect 147644 4508 147700 4564
rect 147308 2604 147364 2660
rect 148652 4732 148708 4788
rect 148092 4450 148148 4452
rect 148092 4398 148094 4450
rect 148094 4398 148146 4450
rect 148146 4398 148148 4450
rect 148092 4396 148148 4398
rect 151340 8428 151396 8484
rect 148988 6748 149044 6804
rect 148764 4508 148820 4564
rect 148204 3836 148260 3892
rect 148092 3612 148148 3668
rect 147980 3276 148036 3332
rect 147756 1260 147812 1316
rect 149548 5852 149604 5908
rect 149100 4508 149156 4564
rect 149100 4338 149156 4340
rect 149100 4286 149102 4338
rect 149102 4286 149154 4338
rect 149154 4286 149156 4338
rect 149100 4284 149156 4286
rect 148652 4060 148708 4116
rect 148876 3724 148932 3780
rect 148316 2492 148372 2548
rect 149324 3612 149380 3668
rect 148988 3554 149044 3556
rect 148988 3502 148990 3554
rect 148990 3502 149042 3554
rect 149042 3502 149044 3554
rect 148988 3500 149044 3502
rect 149660 4450 149716 4452
rect 149660 4398 149662 4450
rect 149662 4398 149714 4450
rect 149714 4398 149716 4450
rect 149660 4396 149716 4398
rect 149772 4284 149828 4340
rect 149772 3948 149828 4004
rect 149772 3612 149828 3668
rect 149996 4844 150052 4900
rect 149996 3724 150052 3780
rect 149884 3388 149940 3444
rect 150668 4898 150724 4900
rect 150668 4846 150670 4898
rect 150670 4846 150722 4898
rect 150722 4846 150724 4898
rect 150668 4844 150724 4846
rect 150556 3836 150612 3892
rect 152572 6524 152628 6580
rect 151004 4284 151060 4340
rect 151452 4338 151508 4340
rect 151452 4286 151454 4338
rect 151454 4286 151506 4338
rect 151506 4286 151508 4338
rect 151452 4284 151508 4286
rect 150444 3500 150500 3556
rect 150780 2940 150836 2996
rect 151676 4172 151732 4228
rect 151116 3948 151172 4004
rect 151116 3724 151172 3780
rect 152012 3724 152068 3780
rect 151900 3554 151956 3556
rect 151900 3502 151902 3554
rect 151902 3502 151954 3554
rect 151954 3502 151956 3554
rect 151900 3500 151956 3502
rect 152124 3388 152180 3444
rect 152460 3388 152516 3444
rect 152796 3612 152852 3668
rect 152684 3500 152740 3556
rect 152908 3442 152964 3444
rect 152908 3390 152910 3442
rect 152910 3390 152962 3442
rect 152962 3390 152964 3442
rect 152908 3388 152964 3390
rect 153692 3554 153748 3556
rect 153692 3502 153694 3554
rect 153694 3502 153746 3554
rect 153746 3502 153748 3554
rect 153692 3500 153748 3502
rect 154028 3500 154084 3556
rect 154364 3612 154420 3668
rect 153916 3388 153972 3444
rect 153468 1148 153524 1204
rect 154588 3388 154644 3444
rect 154700 3330 154756 3332
rect 154700 3278 154702 3330
rect 154702 3278 154754 3330
rect 154754 3278 154756 3330
rect 154700 3276 154756 3278
rect 158076 10218 158132 10220
rect 158076 10166 158078 10218
rect 158078 10166 158130 10218
rect 158130 10166 158132 10218
rect 158076 10164 158132 10166
rect 158180 10218 158236 10220
rect 158180 10166 158182 10218
rect 158182 10166 158234 10218
rect 158234 10166 158236 10218
rect 158180 10164 158236 10166
rect 158284 10218 158340 10220
rect 158284 10166 158286 10218
rect 158286 10166 158338 10218
rect 158338 10166 158340 10218
rect 158284 10164 158340 10166
rect 158076 8650 158132 8652
rect 158076 8598 158078 8650
rect 158078 8598 158130 8650
rect 158130 8598 158132 8650
rect 158076 8596 158132 8598
rect 158180 8650 158236 8652
rect 158180 8598 158182 8650
rect 158182 8598 158234 8650
rect 158234 8598 158236 8650
rect 158180 8596 158236 8598
rect 158284 8650 158340 8652
rect 158284 8598 158286 8650
rect 158286 8598 158338 8650
rect 158338 8598 158340 8650
rect 158284 8596 158340 8598
rect 159068 8092 159124 8148
rect 158076 7082 158132 7084
rect 158076 7030 158078 7082
rect 158078 7030 158130 7082
rect 158130 7030 158132 7082
rect 158076 7028 158132 7030
rect 158180 7082 158236 7084
rect 158180 7030 158182 7082
rect 158182 7030 158234 7082
rect 158234 7030 158236 7082
rect 158180 7028 158236 7030
rect 158284 7082 158340 7084
rect 158284 7030 158286 7082
rect 158286 7030 158338 7082
rect 158338 7030 158340 7082
rect 158284 7028 158340 7030
rect 158076 5514 158132 5516
rect 158076 5462 158078 5514
rect 158078 5462 158130 5514
rect 158130 5462 158132 5514
rect 158076 5460 158132 5462
rect 158180 5514 158236 5516
rect 158180 5462 158182 5514
rect 158182 5462 158234 5514
rect 158234 5462 158236 5514
rect 158180 5460 158236 5462
rect 158284 5514 158340 5516
rect 158284 5462 158286 5514
rect 158286 5462 158338 5514
rect 158338 5462 158340 5514
rect 158284 5460 158340 5462
rect 155372 3612 155428 3668
rect 155820 3612 155876 3668
rect 155484 3500 155540 3556
rect 155036 3442 155092 3444
rect 155036 3390 155038 3442
rect 155038 3390 155090 3442
rect 155090 3390 155092 3442
rect 155036 3388 155092 3390
rect 155596 1484 155652 1540
rect 156492 3836 156548 3892
rect 156716 3554 156772 3556
rect 156716 3502 156718 3554
rect 156718 3502 156770 3554
rect 156770 3502 156772 3554
rect 156716 3500 156772 3502
rect 156604 3388 156660 3444
rect 157164 3388 157220 3444
rect 157388 4396 157444 4452
rect 158076 3946 158132 3948
rect 158076 3894 158078 3946
rect 158078 3894 158130 3946
rect 158130 3894 158132 3946
rect 158076 3892 158132 3894
rect 158180 3946 158236 3948
rect 158180 3894 158182 3946
rect 158182 3894 158234 3946
rect 158234 3894 158236 3946
rect 158180 3892 158236 3894
rect 158284 3946 158340 3948
rect 158284 3894 158286 3946
rect 158286 3894 158338 3946
rect 158338 3894 158340 3946
rect 158284 3892 158340 3894
rect 157724 3500 157780 3556
rect 159516 5628 159572 5684
rect 158508 3500 158564 3556
rect 158956 3554 159012 3556
rect 158956 3502 158958 3554
rect 158958 3502 159010 3554
rect 159010 3502 159012 3554
rect 158956 3500 159012 3502
rect 158844 3388 158900 3444
rect 158620 1372 158676 1428
rect 159292 3388 159348 3444
rect 159404 3500 159460 3556
rect 159180 3276 159236 3332
rect 159852 3442 159908 3444
rect 159852 3390 159854 3442
rect 159854 3390 159906 3442
rect 159906 3390 159908 3442
rect 159852 3388 159908 3390
rect 161420 12012 161476 12068
rect 161084 4284 161140 4340
rect 160636 3554 160692 3556
rect 160636 3502 160638 3554
rect 160638 3502 160690 3554
rect 160690 3502 160692 3554
rect 160636 3500 160692 3502
rect 160524 3388 160580 3444
rect 161532 4338 161588 4340
rect 161532 4286 161534 4338
rect 161534 4286 161586 4338
rect 161586 4286 161588 4338
rect 161532 4284 161588 4286
rect 161644 3388 161700 3444
rect 162764 3500 162820 3556
rect 162204 3388 162260 3444
rect 162540 2268 162596 2324
rect 162876 3442 162932 3444
rect 162876 3390 162878 3442
rect 162878 3390 162930 3442
rect 162930 3390 162932 3442
rect 162876 3388 162932 3390
rect 164332 7532 164388 7588
rect 163660 3554 163716 3556
rect 163660 3502 163662 3554
rect 163662 3502 163714 3554
rect 163714 3502 163716 3554
rect 163660 3500 163716 3502
rect 164108 3500 164164 3556
rect 163884 3388 163940 3444
rect 164444 3500 164500 3556
rect 164668 3442 164724 3444
rect 164668 3390 164670 3442
rect 164670 3390 164722 3442
rect 164722 3390 164724 3442
rect 164668 3388 164724 3390
rect 165452 3554 165508 3556
rect 165452 3502 165454 3554
rect 165454 3502 165506 3554
rect 165506 3502 165508 3554
rect 165452 3500 165508 3502
rect 165788 3500 165844 3556
rect 166124 3500 166180 3556
rect 165676 3388 165732 3444
rect 165228 3330 165284 3332
rect 165228 3278 165230 3330
rect 165230 3278 165282 3330
rect 165282 3278 165284 3330
rect 165228 3276 165284 3278
rect 166348 3388 166404 3444
rect 166460 2380 166516 2436
rect 167132 3500 167188 3556
rect 166796 3442 166852 3444
rect 166796 3390 166798 3442
rect 166798 3390 166850 3442
rect 166850 3390 166852 3442
rect 166796 3388 166852 3390
rect 167244 3388 167300 3444
rect 173436 23546 173492 23548
rect 173436 23494 173438 23546
rect 173438 23494 173490 23546
rect 173490 23494 173492 23546
rect 173436 23492 173492 23494
rect 173540 23546 173596 23548
rect 173540 23494 173542 23546
rect 173542 23494 173594 23546
rect 173594 23494 173596 23546
rect 173540 23492 173596 23494
rect 173644 23546 173700 23548
rect 173644 23494 173646 23546
rect 173646 23494 173698 23546
rect 173698 23494 173700 23546
rect 173644 23492 173700 23494
rect 173436 21978 173492 21980
rect 173436 21926 173438 21978
rect 173438 21926 173490 21978
rect 173490 21926 173492 21978
rect 173436 21924 173492 21926
rect 173540 21978 173596 21980
rect 173540 21926 173542 21978
rect 173542 21926 173594 21978
rect 173594 21926 173596 21978
rect 173540 21924 173596 21926
rect 173644 21978 173700 21980
rect 173644 21926 173646 21978
rect 173646 21926 173698 21978
rect 173698 21926 173700 21978
rect 173644 21924 173700 21926
rect 173436 20410 173492 20412
rect 173436 20358 173438 20410
rect 173438 20358 173490 20410
rect 173490 20358 173492 20410
rect 173436 20356 173492 20358
rect 173540 20410 173596 20412
rect 173540 20358 173542 20410
rect 173542 20358 173594 20410
rect 173594 20358 173596 20410
rect 173540 20356 173596 20358
rect 173644 20410 173700 20412
rect 173644 20358 173646 20410
rect 173646 20358 173698 20410
rect 173698 20358 173700 20410
rect 173644 20356 173700 20358
rect 167804 3612 167860 3668
rect 167580 3554 167636 3556
rect 167580 3502 167582 3554
rect 167582 3502 167634 3554
rect 167634 3502 167636 3554
rect 167580 3500 167636 3502
rect 173436 18842 173492 18844
rect 173436 18790 173438 18842
rect 173438 18790 173490 18842
rect 173490 18790 173492 18842
rect 173436 18788 173492 18790
rect 173540 18842 173596 18844
rect 173540 18790 173542 18842
rect 173542 18790 173594 18842
rect 173594 18790 173596 18842
rect 173540 18788 173596 18790
rect 173644 18842 173700 18844
rect 173644 18790 173646 18842
rect 173646 18790 173698 18842
rect 173698 18790 173700 18842
rect 173644 18788 173700 18790
rect 173436 17274 173492 17276
rect 173436 17222 173438 17274
rect 173438 17222 173490 17274
rect 173490 17222 173492 17274
rect 173436 17220 173492 17222
rect 173540 17274 173596 17276
rect 173540 17222 173542 17274
rect 173542 17222 173594 17274
rect 173594 17222 173596 17274
rect 173540 17220 173596 17222
rect 173644 17274 173700 17276
rect 173644 17222 173646 17274
rect 173646 17222 173698 17274
rect 173698 17222 173700 17274
rect 173644 17220 173700 17222
rect 173436 15706 173492 15708
rect 173436 15654 173438 15706
rect 173438 15654 173490 15706
rect 173490 15654 173492 15706
rect 173436 15652 173492 15654
rect 173540 15706 173596 15708
rect 173540 15654 173542 15706
rect 173542 15654 173594 15706
rect 173594 15654 173596 15706
rect 173540 15652 173596 15654
rect 173644 15706 173700 15708
rect 173644 15654 173646 15706
rect 173646 15654 173698 15706
rect 173698 15654 173700 15706
rect 173644 15652 173700 15654
rect 173436 14138 173492 14140
rect 173436 14086 173438 14138
rect 173438 14086 173490 14138
rect 173490 14086 173492 14138
rect 173436 14084 173492 14086
rect 173540 14138 173596 14140
rect 173540 14086 173542 14138
rect 173542 14086 173594 14138
rect 173594 14086 173596 14138
rect 173540 14084 173596 14086
rect 173644 14138 173700 14140
rect 173644 14086 173646 14138
rect 173646 14086 173698 14138
rect 173698 14086 173700 14138
rect 173644 14084 173700 14086
rect 173436 12570 173492 12572
rect 173436 12518 173438 12570
rect 173438 12518 173490 12570
rect 173490 12518 173492 12570
rect 173436 12516 173492 12518
rect 173540 12570 173596 12572
rect 173540 12518 173542 12570
rect 173542 12518 173594 12570
rect 173594 12518 173596 12570
rect 173540 12516 173596 12518
rect 173644 12570 173700 12572
rect 173644 12518 173646 12570
rect 173646 12518 173698 12570
rect 173698 12518 173700 12570
rect 173644 12516 173700 12518
rect 170380 11900 170436 11956
rect 169260 4844 169316 4900
rect 168140 3388 168196 3444
rect 168588 3442 168644 3444
rect 168588 3390 168590 3442
rect 168590 3390 168642 3442
rect 168642 3390 168644 3442
rect 168588 3388 168644 3390
rect 168252 2716 168308 2772
rect 169260 4396 169316 4452
rect 169036 1596 169092 1652
rect 169484 3612 169540 3668
rect 169596 3500 169652 3556
rect 173436 11002 173492 11004
rect 173436 10950 173438 11002
rect 173438 10950 173490 11002
rect 173490 10950 173492 11002
rect 173436 10948 173492 10950
rect 173540 11002 173596 11004
rect 173540 10950 173542 11002
rect 173542 10950 173594 11002
rect 173594 10950 173596 11002
rect 173540 10948 173596 10950
rect 173644 11002 173700 11004
rect 173644 10950 173646 11002
rect 173646 10950 173698 11002
rect 173698 10950 173700 11002
rect 173644 10948 173700 10950
rect 172172 10332 172228 10388
rect 171276 7980 171332 8036
rect 170716 3554 170772 3556
rect 170716 3502 170718 3554
rect 170718 3502 170770 3554
rect 170770 3502 170772 3554
rect 170716 3500 170772 3502
rect 171164 3500 171220 3556
rect 170604 3388 170660 3444
rect 171388 3388 171444 3444
rect 171612 3442 171668 3444
rect 171612 3390 171614 3442
rect 171614 3390 171666 3442
rect 171666 3390 171668 3442
rect 171612 3388 171668 3390
rect 173436 9434 173492 9436
rect 173436 9382 173438 9434
rect 173438 9382 173490 9434
rect 173490 9382 173492 9434
rect 173436 9380 173492 9382
rect 173540 9434 173596 9436
rect 173540 9382 173542 9434
rect 173542 9382 173594 9434
rect 173594 9382 173596 9434
rect 173540 9380 173596 9382
rect 173644 9434 173700 9436
rect 173644 9382 173646 9434
rect 173646 9382 173698 9434
rect 173698 9382 173700 9434
rect 173644 9380 173700 9382
rect 173436 7866 173492 7868
rect 173436 7814 173438 7866
rect 173438 7814 173490 7866
rect 173490 7814 173492 7866
rect 173436 7812 173492 7814
rect 173540 7866 173596 7868
rect 173540 7814 173542 7866
rect 173542 7814 173594 7866
rect 173594 7814 173596 7866
rect 173540 7812 173596 7814
rect 173644 7866 173700 7868
rect 173644 7814 173646 7866
rect 173646 7814 173698 7866
rect 173698 7814 173700 7866
rect 173644 7812 173700 7814
rect 173436 6298 173492 6300
rect 173436 6246 173438 6298
rect 173438 6246 173490 6298
rect 173490 6246 173492 6298
rect 173436 6244 173492 6246
rect 173540 6298 173596 6300
rect 173540 6246 173542 6298
rect 173542 6246 173594 6298
rect 173594 6246 173596 6298
rect 173540 6244 173596 6246
rect 173644 6298 173700 6300
rect 173644 6246 173646 6298
rect 173646 6246 173698 6298
rect 173698 6246 173700 6298
rect 173644 6244 173700 6246
rect 173180 5292 173236 5348
rect 172396 3554 172452 3556
rect 172396 3502 172398 3554
rect 172398 3502 172450 3554
rect 172450 3502 172452 3554
rect 172396 3500 172452 3502
rect 172284 3388 172340 3444
rect 173436 4730 173492 4732
rect 173436 4678 173438 4730
rect 173438 4678 173490 4730
rect 173490 4678 173492 4730
rect 173436 4676 173492 4678
rect 173540 4730 173596 4732
rect 173540 4678 173542 4730
rect 173542 4678 173594 4730
rect 173594 4678 173596 4730
rect 173540 4676 173596 4678
rect 173644 4730 173700 4732
rect 173644 4678 173646 4730
rect 173646 4678 173698 4730
rect 173698 4678 173700 4730
rect 173644 4676 173700 4678
rect 173404 3388 173460 3444
rect 173964 3276 174020 3332
rect 173436 3162 173492 3164
rect 173436 3110 173438 3162
rect 173438 3110 173490 3162
rect 173490 3110 173492 3162
rect 173436 3108 173492 3110
rect 173540 3162 173596 3164
rect 173540 3110 173542 3162
rect 173542 3110 173594 3162
rect 173594 3110 173596 3162
rect 173540 3108 173596 3110
rect 173644 3162 173700 3164
rect 173644 3110 173646 3162
rect 173646 3110 173698 3162
rect 173698 3110 173700 3162
rect 173644 3108 173700 3110
rect 174972 3330 175028 3332
rect 174972 3278 174974 3330
rect 174974 3278 175026 3330
rect 175026 3278 175028 3330
rect 174972 3276 175028 3278
rect 130508 700 130564 756
<< metal3 >>
rect 26450 117180 26460 117236
rect 26516 117180 27356 117236
rect 27412 117180 27422 117236
rect 49970 117180 49980 117236
rect 50036 117180 50876 117236
rect 50932 117180 50942 117236
rect 144050 117180 144060 117236
rect 144116 117180 144956 117236
rect 145012 117180 145022 117236
rect 167570 117068 167580 117124
rect 167636 117068 168476 117124
rect 168532 117068 168542 117124
rect 4498 116956 4508 117012
rect 4564 116956 5964 117012
rect 6020 116956 6030 117012
rect 54674 116956 54684 117012
rect 54740 116956 55468 117012
rect 55524 116956 55534 117012
rect 153458 116956 153468 117012
rect 153524 116956 155372 117012
rect 155428 116956 155438 117012
rect 4466 116788 4476 116844
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4740 116788 4750 116844
rect 35186 116788 35196 116844
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35460 116788 35470 116844
rect 65906 116788 65916 116844
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 66180 116788 66190 116844
rect 96626 116788 96636 116844
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96900 116788 96910 116844
rect 127346 116788 127356 116844
rect 127412 116788 127460 116844
rect 127516 116788 127564 116844
rect 127620 116788 127630 116844
rect 158066 116788 158076 116844
rect 158132 116788 158180 116844
rect 158236 116788 158284 116844
rect 158340 116788 158350 116844
rect 7634 116620 7644 116676
rect 7700 116620 8428 116676
rect 8484 116620 8494 116676
rect 31154 116620 31164 116676
rect 31220 116620 31948 116676
rect 32004 116620 32014 116676
rect 78194 116620 78204 116676
rect 78260 116620 78988 116676
rect 79044 116620 79054 116676
rect 92306 116620 92316 116676
rect 92372 116620 93212 116676
rect 93268 116620 93278 116676
rect 101714 116620 101724 116676
rect 101780 116620 102508 116676
rect 102564 116620 102574 116676
rect 115826 116620 115836 116676
rect 115892 116620 116732 116676
rect 116788 116620 116798 116676
rect 125234 116620 125244 116676
rect 125300 116620 126028 116676
rect 126084 116620 126094 116676
rect 139346 116620 139356 116676
rect 139412 116620 140252 116676
rect 140308 116620 140318 116676
rect 148754 116620 148764 116676
rect 148820 116620 149548 116676
rect 149604 116620 149614 116676
rect 162866 116620 162876 116676
rect 162932 116620 163772 116676
rect 163828 116620 163838 116676
rect 172274 116620 172284 116676
rect 172340 116620 173068 116676
rect 173124 116620 173134 116676
rect 2930 116508 2940 116564
rect 2996 116508 3388 116564
rect 3444 116508 3454 116564
rect 9202 116508 9212 116564
rect 9268 116508 10108 116564
rect 10164 116508 10174 116564
rect 28018 116508 28028 116564
rect 28084 116508 29484 116564
rect 29540 116508 29550 116564
rect 32722 116508 32732 116564
rect 32788 116508 33628 116564
rect 33684 116508 33694 116564
rect 51538 116508 51548 116564
rect 51604 116508 53004 116564
rect 53060 116508 53070 116564
rect 56242 116508 56252 116564
rect 56308 116508 57148 116564
rect 57204 116508 57214 116564
rect 67172 116508 73052 116564
rect 73108 116508 73118 116564
rect 73490 116508 73500 116564
rect 73556 116508 74396 116564
rect 74452 116508 74462 116564
rect 75058 116508 75068 116564
rect 75124 116508 76524 116564
rect 76580 116508 76590 116564
rect 79762 116508 79772 116564
rect 79828 116508 80668 116564
rect 80724 116508 80734 116564
rect 97010 116508 97020 116564
rect 97076 116508 97916 116564
rect 97972 116508 97982 116564
rect 98578 116508 98588 116564
rect 98644 116508 100044 116564
rect 100100 116508 100110 116564
rect 103282 116508 103292 116564
rect 103348 116508 104188 116564
rect 104244 116508 104254 116564
rect 106418 116508 106428 116564
rect 106484 116508 108332 116564
rect 108388 116508 108398 116564
rect 120530 116508 120540 116564
rect 120596 116508 121436 116564
rect 121492 116508 121502 116564
rect 122098 116508 122108 116564
rect 122164 116508 124012 116564
rect 124068 116508 124078 116564
rect 126802 116508 126812 116564
rect 126868 116508 127932 116564
rect 127988 116508 127998 116564
rect 129938 116508 129948 116564
rect 130004 116508 131852 116564
rect 131908 116508 131918 116564
rect 145618 116508 145628 116564
rect 145684 116508 147532 116564
rect 147588 116508 147598 116564
rect 150322 116508 150332 116564
rect 150388 116508 151452 116564
rect 151508 116508 151518 116564
rect 18050 116396 18060 116452
rect 18116 116396 19852 116452
rect 19908 116396 20524 116452
rect 20580 116396 20590 116452
rect 48066 116396 48076 116452
rect 48132 116396 48748 116452
rect 48804 116396 48814 116452
rect 67172 116340 67228 116508
rect 106306 116396 106316 116452
rect 106372 116396 107660 116452
rect 107716 116396 107726 116452
rect 120082 116396 120092 116452
rect 120148 116396 126028 116452
rect 129826 116396 129836 116452
rect 129892 116396 131180 116452
rect 131236 116396 131246 116452
rect 137732 116396 146076 116452
rect 146132 116396 146860 116452
rect 146916 116396 146926 116452
rect 153458 116396 153468 116452
rect 153524 116396 154700 116452
rect 154756 116396 154766 116452
rect 170930 116396 170940 116452
rect 170996 116396 172284 116452
rect 172340 116396 172350 116452
rect 38882 116284 38892 116340
rect 38948 116284 39340 116340
rect 39396 116284 67228 116340
rect 125972 116340 126028 116396
rect 137732 116340 137788 116396
rect 125972 116284 137788 116340
rect 164434 116284 164444 116340
rect 164500 116284 164892 116340
rect 164948 116284 164958 116340
rect 169138 116284 169148 116340
rect 169204 116284 170380 116340
rect 170436 116284 170446 116340
rect 10882 116172 10892 116228
rect 10948 116172 11340 116228
rect 11396 116172 12684 116228
rect 12740 116172 12750 116228
rect 67106 116172 67116 116228
rect 67172 116172 67564 116228
rect 67620 116172 69916 116228
rect 69972 116172 69982 116228
rect 71362 116172 71372 116228
rect 71428 116172 72268 116228
rect 72324 116172 72334 116228
rect 90626 116172 90636 116228
rect 90692 116172 91084 116228
rect 91140 116172 95340 116228
rect 95396 116172 95406 116228
rect 104962 116172 104972 116228
rect 105028 116172 105420 116228
rect 105476 116172 106092 116228
rect 106148 116172 106158 116228
rect 118962 116172 118972 116228
rect 119028 116172 122556 116228
rect 122612 116172 123340 116228
rect 123396 116172 123406 116228
rect 57922 116060 57932 116116
rect 57988 116060 58380 116116
rect 58436 116060 80220 116116
rect 80276 116060 80286 116116
rect 85922 116060 85932 116116
rect 85988 116060 86380 116116
rect 86436 116060 90860 116116
rect 90916 116060 90926 116116
rect 19826 116004 19836 116060
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 20100 116004 20110 116060
rect 50546 116004 50556 116060
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50820 116004 50830 116060
rect 81266 116004 81276 116060
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81540 116004 81550 116060
rect 111986 116004 111996 116060
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 112260 116004 112270 116060
rect 142706 116004 142716 116060
rect 142772 116004 142820 116060
rect 142876 116004 142924 116060
rect 142980 116004 142990 116060
rect 173426 116004 173436 116060
rect 173492 116004 173540 116060
rect 173596 116004 173644 116060
rect 173700 116004 173710 116060
rect 12338 115836 12348 115892
rect 12404 115836 13244 115892
rect 13300 115836 13310 115892
rect 17042 115836 17052 115892
rect 17108 115836 18620 115892
rect 18676 115836 18686 115892
rect 35858 115836 35868 115892
rect 35924 115836 36764 115892
rect 36820 115836 36830 115892
rect 40674 115836 40684 115892
rect 40740 115836 42252 115892
rect 42308 115836 42318 115892
rect 59378 115836 59388 115892
rect 59444 115836 60284 115892
rect 60340 115836 60350 115892
rect 82898 115836 82908 115892
rect 82964 115836 83804 115892
rect 83860 115836 83870 115892
rect 178098 115836 178108 115892
rect 178164 115836 178556 115892
rect 178612 115836 178622 115892
rect 53778 115724 53788 115780
rect 53844 115724 55132 115780
rect 55188 115724 55198 115780
rect 93874 115724 93884 115780
rect 93940 115724 94444 115780
rect 94500 115724 94510 115780
rect 107986 115724 107996 115780
rect 108052 115724 108556 115780
rect 108612 115724 108622 115780
rect 117394 115724 117404 115780
rect 117460 115724 118524 115780
rect 118580 115724 118590 115780
rect 131506 115724 131516 115780
rect 131572 115724 132636 115780
rect 132692 115724 132702 115780
rect 140914 115724 140924 115780
rect 140980 115724 142044 115780
rect 142100 115724 142110 115780
rect 5170 115612 5180 115668
rect 5236 115612 7196 115668
rect 7252 115612 7980 115668
rect 8036 115612 11116 115668
rect 11172 115612 11676 115668
rect 11732 115612 16044 115668
rect 16100 115612 16716 115668
rect 16772 115612 20860 115668
rect 20916 115612 21532 115668
rect 21588 115612 25564 115668
rect 25620 115612 26236 115668
rect 26292 115612 30268 115668
rect 30324 115612 30940 115668
rect 30996 115612 34636 115668
rect 34692 115612 35196 115668
rect 35252 115612 39676 115668
rect 39732 115612 40236 115668
rect 40292 115612 44380 115668
rect 44436 115612 45052 115668
rect 45108 115612 48748 115668
rect 48804 115612 49756 115668
rect 49812 115612 54460 115668
rect 54516 115612 58212 115668
rect 91410 115612 91420 115668
rect 91476 115612 91980 115668
rect 92036 115612 96460 115668
rect 96516 115612 97580 115668
rect 97636 115612 100828 115668
rect 100884 115612 101388 115668
rect 101444 115612 105420 115668
rect 105476 115612 105980 115668
rect 106036 115612 110460 115668
rect 110516 115612 110796 115668
rect 110852 115612 114940 115668
rect 114996 115612 115500 115668
rect 115556 115612 120316 115668
rect 120372 115612 121324 115668
rect 121380 115612 124236 115668
rect 124292 115612 124796 115668
rect 124852 115612 128940 115668
rect 128996 115612 129612 115668
rect 129668 115612 133756 115668
rect 133812 115612 134316 115668
rect 134372 115612 138460 115668
rect 138516 115612 139132 115668
rect 139188 115612 143164 115668
rect 143220 115612 143836 115668
rect 143892 115612 147868 115668
rect 147924 115612 148540 115668
rect 148596 115612 152124 115668
rect 152180 115612 153244 115668
rect 153300 115612 157276 115668
rect 157332 115612 157836 115668
rect 157892 115612 161980 115668
rect 162036 115612 162540 115668
rect 162596 115612 166684 115668
rect 166740 115612 167244 115668
rect 167300 115612 170044 115668
rect 170100 115612 170604 115668
rect 170660 115612 170670 115668
rect 53788 115556 53844 115612
rect 58156 115556 58212 115612
rect 53778 115500 53788 115556
rect 53844 115500 53854 115556
rect 58146 115500 58156 115556
rect 58212 115500 58716 115556
rect 58772 115500 63196 115556
rect 63252 115500 63756 115556
rect 63812 115500 67900 115556
rect 67956 115500 68572 115556
rect 68628 115500 72604 115556
rect 72660 115500 73500 115556
rect 73556 115500 77308 115556
rect 77364 115500 77980 115556
rect 78036 115500 81676 115556
rect 81732 115500 82236 115556
rect 82292 115500 82302 115556
rect 95330 115500 95340 115556
rect 95396 115500 95900 115556
rect 95956 115500 97468 115556
rect 97524 115500 97534 115556
rect 113026 115500 113036 115556
rect 113092 115500 113932 115556
rect 113988 115500 114380 115556
rect 114436 115500 114446 115556
rect 125234 115500 125244 115556
rect 125300 115500 126924 115556
rect 126980 115500 126990 115556
rect 4466 115220 4476 115276
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4740 115220 4750 115276
rect 35186 115220 35196 115276
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35460 115220 35470 115276
rect 65906 115220 65916 115276
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 66180 115220 66190 115276
rect 96626 115220 96636 115276
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96900 115220 96910 115276
rect 127346 115220 127356 115276
rect 127412 115220 127460 115276
rect 127516 115220 127564 115276
rect 127620 115220 127630 115276
rect 158066 115220 158076 115276
rect 158132 115220 158180 115276
rect 158236 115220 158284 115276
rect 158340 115220 158350 115276
rect 64194 115052 64204 115108
rect 64260 115052 64988 115108
rect 65044 115052 65054 115108
rect 82226 114828 82236 114884
rect 82292 114828 86716 114884
rect 86772 114828 87612 114884
rect 87668 114828 91420 114884
rect 91476 114828 91486 114884
rect 19826 114436 19836 114492
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 20100 114436 20110 114492
rect 50546 114436 50556 114492
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50820 114436 50830 114492
rect 81266 114436 81276 114492
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81540 114436 81550 114492
rect 111986 114436 111996 114492
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 112260 114436 112270 114492
rect 142706 114436 142716 114492
rect 142772 114436 142820 114492
rect 142876 114436 142924 114492
rect 142980 114436 142990 114492
rect 173426 114436 173436 114492
rect 173492 114436 173540 114492
rect 173596 114436 173644 114492
rect 173700 114436 173710 114492
rect 4466 113652 4476 113708
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4740 113652 4750 113708
rect 35186 113652 35196 113708
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35460 113652 35470 113708
rect 65906 113652 65916 113708
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 66180 113652 66190 113708
rect 96626 113652 96636 113708
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96900 113652 96910 113708
rect 127346 113652 127356 113708
rect 127412 113652 127460 113708
rect 127516 113652 127564 113708
rect 127620 113652 127630 113708
rect 158066 113652 158076 113708
rect 158132 113652 158180 113708
rect 158236 113652 158284 113708
rect 158340 113652 158350 113708
rect 19826 112868 19836 112924
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 20100 112868 20110 112924
rect 50546 112868 50556 112924
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50820 112868 50830 112924
rect 81266 112868 81276 112924
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81540 112868 81550 112924
rect 111986 112868 111996 112924
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 112260 112868 112270 112924
rect 142706 112868 142716 112924
rect 142772 112868 142820 112924
rect 142876 112868 142924 112924
rect 142980 112868 142990 112924
rect 173426 112868 173436 112924
rect 173492 112868 173540 112924
rect 173596 112868 173644 112924
rect 173700 112868 173710 112924
rect 4466 112084 4476 112140
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4740 112084 4750 112140
rect 35186 112084 35196 112140
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35460 112084 35470 112140
rect 65906 112084 65916 112140
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 66180 112084 66190 112140
rect 96626 112084 96636 112140
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96900 112084 96910 112140
rect 127346 112084 127356 112140
rect 127412 112084 127460 112140
rect 127516 112084 127564 112140
rect 127620 112084 127630 112140
rect 158066 112084 158076 112140
rect 158132 112084 158180 112140
rect 158236 112084 158284 112140
rect 158340 112084 158350 112140
rect 19826 111300 19836 111356
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 20100 111300 20110 111356
rect 50546 111300 50556 111356
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50820 111300 50830 111356
rect 81266 111300 81276 111356
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81540 111300 81550 111356
rect 111986 111300 111996 111356
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 112260 111300 112270 111356
rect 142706 111300 142716 111356
rect 142772 111300 142820 111356
rect 142876 111300 142924 111356
rect 142980 111300 142990 111356
rect 173426 111300 173436 111356
rect 173492 111300 173540 111356
rect 173596 111300 173644 111356
rect 173700 111300 173710 111356
rect 4466 110516 4476 110572
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4740 110516 4750 110572
rect 35186 110516 35196 110572
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35460 110516 35470 110572
rect 65906 110516 65916 110572
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 66180 110516 66190 110572
rect 96626 110516 96636 110572
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96900 110516 96910 110572
rect 127346 110516 127356 110572
rect 127412 110516 127460 110572
rect 127516 110516 127564 110572
rect 127620 110516 127630 110572
rect 158066 110516 158076 110572
rect 158132 110516 158180 110572
rect 158236 110516 158284 110572
rect 158340 110516 158350 110572
rect 19826 109732 19836 109788
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 20100 109732 20110 109788
rect 50546 109732 50556 109788
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50820 109732 50830 109788
rect 81266 109732 81276 109788
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81540 109732 81550 109788
rect 111986 109732 111996 109788
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 112260 109732 112270 109788
rect 142706 109732 142716 109788
rect 142772 109732 142820 109788
rect 142876 109732 142924 109788
rect 142980 109732 142990 109788
rect 173426 109732 173436 109788
rect 173492 109732 173540 109788
rect 173596 109732 173644 109788
rect 173700 109732 173710 109788
rect 4466 108948 4476 109004
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4740 108948 4750 109004
rect 35186 108948 35196 109004
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35460 108948 35470 109004
rect 65906 108948 65916 109004
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 66180 108948 66190 109004
rect 96626 108948 96636 109004
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96900 108948 96910 109004
rect 127346 108948 127356 109004
rect 127412 108948 127460 109004
rect 127516 108948 127564 109004
rect 127620 108948 127630 109004
rect 158066 108948 158076 109004
rect 158132 108948 158180 109004
rect 158236 108948 158284 109004
rect 158340 108948 158350 109004
rect 6626 108332 6636 108388
rect 6692 108332 57148 108388
rect 57204 108332 57214 108388
rect 19826 108164 19836 108220
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 20100 108164 20110 108220
rect 50546 108164 50556 108220
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50820 108164 50830 108220
rect 81266 108164 81276 108220
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81540 108164 81550 108220
rect 111986 108164 111996 108220
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 112260 108164 112270 108220
rect 142706 108164 142716 108220
rect 142772 108164 142820 108220
rect 142876 108164 142924 108220
rect 142980 108164 142990 108220
rect 173426 108164 173436 108220
rect 173492 108164 173540 108220
rect 173596 108164 173644 108220
rect 173700 108164 173710 108220
rect 4466 107380 4476 107436
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4740 107380 4750 107436
rect 35186 107380 35196 107436
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35460 107380 35470 107436
rect 65906 107380 65916 107436
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 66180 107380 66190 107436
rect 96626 107380 96636 107436
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96900 107380 96910 107436
rect 127346 107380 127356 107436
rect 127412 107380 127460 107436
rect 127516 107380 127564 107436
rect 127620 107380 127630 107436
rect 158066 107380 158076 107436
rect 158132 107380 158180 107436
rect 158236 107380 158284 107436
rect 158340 107380 158350 107436
rect 19826 106596 19836 106652
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 20100 106596 20110 106652
rect 50546 106596 50556 106652
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50820 106596 50830 106652
rect 81266 106596 81276 106652
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81540 106596 81550 106652
rect 111986 106596 111996 106652
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 112260 106596 112270 106652
rect 142706 106596 142716 106652
rect 142772 106596 142820 106652
rect 142876 106596 142924 106652
rect 142980 106596 142990 106652
rect 173426 106596 173436 106652
rect 173492 106596 173540 106652
rect 173596 106596 173644 106652
rect 173700 106596 173710 106652
rect 4466 105812 4476 105868
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4740 105812 4750 105868
rect 35186 105812 35196 105868
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35460 105812 35470 105868
rect 65906 105812 65916 105868
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 66180 105812 66190 105868
rect 96626 105812 96636 105868
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96900 105812 96910 105868
rect 127346 105812 127356 105868
rect 127412 105812 127460 105868
rect 127516 105812 127564 105868
rect 127620 105812 127630 105868
rect 158066 105812 158076 105868
rect 158132 105812 158180 105868
rect 158236 105812 158284 105868
rect 158340 105812 158350 105868
rect 19826 105028 19836 105084
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 20100 105028 20110 105084
rect 50546 105028 50556 105084
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50820 105028 50830 105084
rect 81266 105028 81276 105084
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81540 105028 81550 105084
rect 111986 105028 111996 105084
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 112260 105028 112270 105084
rect 142706 105028 142716 105084
rect 142772 105028 142820 105084
rect 142876 105028 142924 105084
rect 142980 105028 142990 105084
rect 173426 105028 173436 105084
rect 173492 105028 173540 105084
rect 173596 105028 173644 105084
rect 173700 105028 173710 105084
rect 4466 104244 4476 104300
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4740 104244 4750 104300
rect 35186 104244 35196 104300
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35460 104244 35470 104300
rect 65906 104244 65916 104300
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 66180 104244 66190 104300
rect 96626 104244 96636 104300
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96900 104244 96910 104300
rect 127346 104244 127356 104300
rect 127412 104244 127460 104300
rect 127516 104244 127564 104300
rect 127620 104244 127630 104300
rect 158066 104244 158076 104300
rect 158132 104244 158180 104300
rect 158236 104244 158284 104300
rect 158340 104244 158350 104300
rect 19826 103460 19836 103516
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 20100 103460 20110 103516
rect 50546 103460 50556 103516
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50820 103460 50830 103516
rect 81266 103460 81276 103516
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81540 103460 81550 103516
rect 111986 103460 111996 103516
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 112260 103460 112270 103516
rect 142706 103460 142716 103516
rect 142772 103460 142820 103516
rect 142876 103460 142924 103516
rect 142980 103460 142990 103516
rect 173426 103460 173436 103516
rect 173492 103460 173540 103516
rect 173596 103460 173644 103516
rect 173700 103460 173710 103516
rect 4466 102676 4476 102732
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4740 102676 4750 102732
rect 35186 102676 35196 102732
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35460 102676 35470 102732
rect 65906 102676 65916 102732
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 66180 102676 66190 102732
rect 96626 102676 96636 102732
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96900 102676 96910 102732
rect 127346 102676 127356 102732
rect 127412 102676 127460 102732
rect 127516 102676 127564 102732
rect 127620 102676 127630 102732
rect 158066 102676 158076 102732
rect 158132 102676 158180 102732
rect 158236 102676 158284 102732
rect 158340 102676 158350 102732
rect 19826 101892 19836 101948
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 20100 101892 20110 101948
rect 50546 101892 50556 101948
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50820 101892 50830 101948
rect 81266 101892 81276 101948
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81540 101892 81550 101948
rect 111986 101892 111996 101948
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 112260 101892 112270 101948
rect 142706 101892 142716 101948
rect 142772 101892 142820 101948
rect 142876 101892 142924 101948
rect 142980 101892 142990 101948
rect 173426 101892 173436 101948
rect 173492 101892 173540 101948
rect 173596 101892 173644 101948
rect 173700 101892 173710 101948
rect 4466 101108 4476 101164
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4740 101108 4750 101164
rect 35186 101108 35196 101164
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35460 101108 35470 101164
rect 65906 101108 65916 101164
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 66180 101108 66190 101164
rect 96626 101108 96636 101164
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96900 101108 96910 101164
rect 127346 101108 127356 101164
rect 127412 101108 127460 101164
rect 127516 101108 127564 101164
rect 127620 101108 127630 101164
rect 158066 101108 158076 101164
rect 158132 101108 158180 101164
rect 158236 101108 158284 101164
rect 158340 101108 158350 101164
rect 19826 100324 19836 100380
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 20100 100324 20110 100380
rect 50546 100324 50556 100380
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50820 100324 50830 100380
rect 81266 100324 81276 100380
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81540 100324 81550 100380
rect 111986 100324 111996 100380
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 112260 100324 112270 100380
rect 142706 100324 142716 100380
rect 142772 100324 142820 100380
rect 142876 100324 142924 100380
rect 142980 100324 142990 100380
rect 173426 100324 173436 100380
rect 173492 100324 173540 100380
rect 173596 100324 173644 100380
rect 173700 100324 173710 100380
rect 4466 99540 4476 99596
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4740 99540 4750 99596
rect 35186 99540 35196 99596
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35460 99540 35470 99596
rect 65906 99540 65916 99596
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 66180 99540 66190 99596
rect 96626 99540 96636 99596
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96900 99540 96910 99596
rect 127346 99540 127356 99596
rect 127412 99540 127460 99596
rect 127516 99540 127564 99596
rect 127620 99540 127630 99596
rect 158066 99540 158076 99596
rect 158132 99540 158180 99596
rect 158236 99540 158284 99596
rect 158340 99540 158350 99596
rect 19826 98756 19836 98812
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 20100 98756 20110 98812
rect 50546 98756 50556 98812
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50820 98756 50830 98812
rect 81266 98756 81276 98812
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81540 98756 81550 98812
rect 111986 98756 111996 98812
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 112260 98756 112270 98812
rect 142706 98756 142716 98812
rect 142772 98756 142820 98812
rect 142876 98756 142924 98812
rect 142980 98756 142990 98812
rect 173426 98756 173436 98812
rect 173492 98756 173540 98812
rect 173596 98756 173644 98812
rect 173700 98756 173710 98812
rect 4466 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4750 98028
rect 35186 97972 35196 98028
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35460 97972 35470 98028
rect 65906 97972 65916 98028
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 66180 97972 66190 98028
rect 96626 97972 96636 98028
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96900 97972 96910 98028
rect 127346 97972 127356 98028
rect 127412 97972 127460 98028
rect 127516 97972 127564 98028
rect 127620 97972 127630 98028
rect 158066 97972 158076 98028
rect 158132 97972 158180 98028
rect 158236 97972 158284 98028
rect 158340 97972 158350 98028
rect 19826 97188 19836 97244
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 20100 97188 20110 97244
rect 50546 97188 50556 97244
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50820 97188 50830 97244
rect 81266 97188 81276 97244
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81540 97188 81550 97244
rect 111986 97188 111996 97244
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 112260 97188 112270 97244
rect 142706 97188 142716 97244
rect 142772 97188 142820 97244
rect 142876 97188 142924 97244
rect 142980 97188 142990 97244
rect 173426 97188 173436 97244
rect 173492 97188 173540 97244
rect 173596 97188 173644 97244
rect 173700 97188 173710 97244
rect 4466 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4750 96460
rect 35186 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35470 96460
rect 65906 96404 65916 96460
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 66180 96404 66190 96460
rect 96626 96404 96636 96460
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96900 96404 96910 96460
rect 127346 96404 127356 96460
rect 127412 96404 127460 96460
rect 127516 96404 127564 96460
rect 127620 96404 127630 96460
rect 158066 96404 158076 96460
rect 158132 96404 158180 96460
rect 158236 96404 158284 96460
rect 158340 96404 158350 96460
rect 19826 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20110 95676
rect 50546 95620 50556 95676
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50820 95620 50830 95676
rect 81266 95620 81276 95676
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81540 95620 81550 95676
rect 111986 95620 111996 95676
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 112260 95620 112270 95676
rect 142706 95620 142716 95676
rect 142772 95620 142820 95676
rect 142876 95620 142924 95676
rect 142980 95620 142990 95676
rect 173426 95620 173436 95676
rect 173492 95620 173540 95676
rect 173596 95620 173644 95676
rect 173700 95620 173710 95676
rect 4466 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4750 94892
rect 35186 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35470 94892
rect 65906 94836 65916 94892
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 66180 94836 66190 94892
rect 96626 94836 96636 94892
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96900 94836 96910 94892
rect 127346 94836 127356 94892
rect 127412 94836 127460 94892
rect 127516 94836 127564 94892
rect 127620 94836 127630 94892
rect 158066 94836 158076 94892
rect 158132 94836 158180 94892
rect 158236 94836 158284 94892
rect 158340 94836 158350 94892
rect 19826 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20110 94108
rect 50546 94052 50556 94108
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50820 94052 50830 94108
rect 81266 94052 81276 94108
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81540 94052 81550 94108
rect 111986 94052 111996 94108
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 112260 94052 112270 94108
rect 142706 94052 142716 94108
rect 142772 94052 142820 94108
rect 142876 94052 142924 94108
rect 142980 94052 142990 94108
rect 173426 94052 173436 94108
rect 173492 94052 173540 94108
rect 173596 94052 173644 94108
rect 173700 94052 173710 94108
rect 4466 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4750 93324
rect 35186 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35470 93324
rect 65906 93268 65916 93324
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 66180 93268 66190 93324
rect 96626 93268 96636 93324
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96900 93268 96910 93324
rect 127346 93268 127356 93324
rect 127412 93268 127460 93324
rect 127516 93268 127564 93324
rect 127620 93268 127630 93324
rect 158066 93268 158076 93324
rect 158132 93268 158180 93324
rect 158236 93268 158284 93324
rect 158340 93268 158350 93324
rect 19826 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20110 92540
rect 50546 92484 50556 92540
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50820 92484 50830 92540
rect 81266 92484 81276 92540
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81540 92484 81550 92540
rect 111986 92484 111996 92540
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 112260 92484 112270 92540
rect 142706 92484 142716 92540
rect 142772 92484 142820 92540
rect 142876 92484 142924 92540
rect 142980 92484 142990 92540
rect 173426 92484 173436 92540
rect 173492 92484 173540 92540
rect 173596 92484 173644 92540
rect 173700 92484 173710 92540
rect 4466 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4750 91756
rect 35186 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35470 91756
rect 65906 91700 65916 91756
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 66180 91700 66190 91756
rect 96626 91700 96636 91756
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96900 91700 96910 91756
rect 127346 91700 127356 91756
rect 127412 91700 127460 91756
rect 127516 91700 127564 91756
rect 127620 91700 127630 91756
rect 158066 91700 158076 91756
rect 158132 91700 158180 91756
rect 158236 91700 158284 91756
rect 158340 91700 158350 91756
rect 19826 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20110 90972
rect 50546 90916 50556 90972
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50820 90916 50830 90972
rect 81266 90916 81276 90972
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81540 90916 81550 90972
rect 111986 90916 111996 90972
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 112260 90916 112270 90972
rect 142706 90916 142716 90972
rect 142772 90916 142820 90972
rect 142876 90916 142924 90972
rect 142980 90916 142990 90972
rect 173426 90916 173436 90972
rect 173492 90916 173540 90972
rect 173596 90916 173644 90972
rect 173700 90916 173710 90972
rect 4466 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4750 90188
rect 35186 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35470 90188
rect 65906 90132 65916 90188
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 66180 90132 66190 90188
rect 96626 90132 96636 90188
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96900 90132 96910 90188
rect 127346 90132 127356 90188
rect 127412 90132 127460 90188
rect 127516 90132 127564 90188
rect 127620 90132 127630 90188
rect 158066 90132 158076 90188
rect 158132 90132 158180 90188
rect 158236 90132 158284 90188
rect 158340 90132 158350 90188
rect 19826 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20110 89404
rect 50546 89348 50556 89404
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50820 89348 50830 89404
rect 81266 89348 81276 89404
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81540 89348 81550 89404
rect 111986 89348 111996 89404
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 112260 89348 112270 89404
rect 142706 89348 142716 89404
rect 142772 89348 142820 89404
rect 142876 89348 142924 89404
rect 142980 89348 142990 89404
rect 173426 89348 173436 89404
rect 173492 89348 173540 89404
rect 173596 89348 173644 89404
rect 173700 89348 173710 89404
rect 4466 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4750 88620
rect 35186 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35470 88620
rect 65906 88564 65916 88620
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 66180 88564 66190 88620
rect 96626 88564 96636 88620
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96900 88564 96910 88620
rect 127346 88564 127356 88620
rect 127412 88564 127460 88620
rect 127516 88564 127564 88620
rect 127620 88564 127630 88620
rect 158066 88564 158076 88620
rect 158132 88564 158180 88620
rect 158236 88564 158284 88620
rect 158340 88564 158350 88620
rect 19826 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20110 87836
rect 50546 87780 50556 87836
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50820 87780 50830 87836
rect 81266 87780 81276 87836
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81540 87780 81550 87836
rect 111986 87780 111996 87836
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 112260 87780 112270 87836
rect 142706 87780 142716 87836
rect 142772 87780 142820 87836
rect 142876 87780 142924 87836
rect 142980 87780 142990 87836
rect 173426 87780 173436 87836
rect 173492 87780 173540 87836
rect 173596 87780 173644 87836
rect 173700 87780 173710 87836
rect 4466 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4750 87052
rect 35186 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35470 87052
rect 65906 86996 65916 87052
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 66180 86996 66190 87052
rect 96626 86996 96636 87052
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96900 86996 96910 87052
rect 127346 86996 127356 87052
rect 127412 86996 127460 87052
rect 127516 86996 127564 87052
rect 127620 86996 127630 87052
rect 158066 86996 158076 87052
rect 158132 86996 158180 87052
rect 158236 86996 158284 87052
rect 158340 86996 158350 87052
rect 19826 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20110 86268
rect 50546 86212 50556 86268
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50820 86212 50830 86268
rect 81266 86212 81276 86268
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81540 86212 81550 86268
rect 111986 86212 111996 86268
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 112260 86212 112270 86268
rect 142706 86212 142716 86268
rect 142772 86212 142820 86268
rect 142876 86212 142924 86268
rect 142980 86212 142990 86268
rect 173426 86212 173436 86268
rect 173492 86212 173540 86268
rect 173596 86212 173644 86268
rect 173700 86212 173710 86268
rect 4466 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4750 85484
rect 35186 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35470 85484
rect 65906 85428 65916 85484
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 66180 85428 66190 85484
rect 96626 85428 96636 85484
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96900 85428 96910 85484
rect 127346 85428 127356 85484
rect 127412 85428 127460 85484
rect 127516 85428 127564 85484
rect 127620 85428 127630 85484
rect 158066 85428 158076 85484
rect 158132 85428 158180 85484
rect 158236 85428 158284 85484
rect 158340 85428 158350 85484
rect 19826 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20110 84700
rect 50546 84644 50556 84700
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50820 84644 50830 84700
rect 81266 84644 81276 84700
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81540 84644 81550 84700
rect 111986 84644 111996 84700
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 112260 84644 112270 84700
rect 142706 84644 142716 84700
rect 142772 84644 142820 84700
rect 142876 84644 142924 84700
rect 142980 84644 142990 84700
rect 173426 84644 173436 84700
rect 173492 84644 173540 84700
rect 173596 84644 173644 84700
rect 173700 84644 173710 84700
rect 4466 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4750 83916
rect 35186 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35470 83916
rect 65906 83860 65916 83916
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 66180 83860 66190 83916
rect 96626 83860 96636 83916
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96900 83860 96910 83916
rect 127346 83860 127356 83916
rect 127412 83860 127460 83916
rect 127516 83860 127564 83916
rect 127620 83860 127630 83916
rect 158066 83860 158076 83916
rect 158132 83860 158180 83916
rect 158236 83860 158284 83916
rect 158340 83860 158350 83916
rect 19826 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20110 83132
rect 50546 83076 50556 83132
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50820 83076 50830 83132
rect 81266 83076 81276 83132
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81540 83076 81550 83132
rect 111986 83076 111996 83132
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 112260 83076 112270 83132
rect 142706 83076 142716 83132
rect 142772 83076 142820 83132
rect 142876 83076 142924 83132
rect 142980 83076 142990 83132
rect 173426 83076 173436 83132
rect 173492 83076 173540 83132
rect 173596 83076 173644 83132
rect 173700 83076 173710 83132
rect 4466 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4750 82348
rect 35186 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35470 82348
rect 65906 82292 65916 82348
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 66180 82292 66190 82348
rect 96626 82292 96636 82348
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96900 82292 96910 82348
rect 127346 82292 127356 82348
rect 127412 82292 127460 82348
rect 127516 82292 127564 82348
rect 127620 82292 127630 82348
rect 158066 82292 158076 82348
rect 158132 82292 158180 82348
rect 158236 82292 158284 82348
rect 158340 82292 158350 82348
rect 19826 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20110 81564
rect 50546 81508 50556 81564
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50820 81508 50830 81564
rect 81266 81508 81276 81564
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81540 81508 81550 81564
rect 111986 81508 111996 81564
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 112260 81508 112270 81564
rect 142706 81508 142716 81564
rect 142772 81508 142820 81564
rect 142876 81508 142924 81564
rect 142980 81508 142990 81564
rect 173426 81508 173436 81564
rect 173492 81508 173540 81564
rect 173596 81508 173644 81564
rect 173700 81508 173710 81564
rect 4466 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4750 80780
rect 35186 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35470 80780
rect 65906 80724 65916 80780
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 66180 80724 66190 80780
rect 96626 80724 96636 80780
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96900 80724 96910 80780
rect 127346 80724 127356 80780
rect 127412 80724 127460 80780
rect 127516 80724 127564 80780
rect 127620 80724 127630 80780
rect 158066 80724 158076 80780
rect 158132 80724 158180 80780
rect 158236 80724 158284 80780
rect 158340 80724 158350 80780
rect 19826 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20110 79996
rect 50546 79940 50556 79996
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50820 79940 50830 79996
rect 81266 79940 81276 79996
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81540 79940 81550 79996
rect 111986 79940 111996 79996
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 112260 79940 112270 79996
rect 142706 79940 142716 79996
rect 142772 79940 142820 79996
rect 142876 79940 142924 79996
rect 142980 79940 142990 79996
rect 173426 79940 173436 79996
rect 173492 79940 173540 79996
rect 173596 79940 173644 79996
rect 173700 79940 173710 79996
rect 4466 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4750 79212
rect 35186 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35470 79212
rect 65906 79156 65916 79212
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 66180 79156 66190 79212
rect 96626 79156 96636 79212
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96900 79156 96910 79212
rect 127346 79156 127356 79212
rect 127412 79156 127460 79212
rect 127516 79156 127564 79212
rect 127620 79156 127630 79212
rect 158066 79156 158076 79212
rect 158132 79156 158180 79212
rect 158236 79156 158284 79212
rect 158340 79156 158350 79212
rect 19826 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20110 78428
rect 50546 78372 50556 78428
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50820 78372 50830 78428
rect 81266 78372 81276 78428
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81540 78372 81550 78428
rect 111986 78372 111996 78428
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 112260 78372 112270 78428
rect 142706 78372 142716 78428
rect 142772 78372 142820 78428
rect 142876 78372 142924 78428
rect 142980 78372 142990 78428
rect 173426 78372 173436 78428
rect 173492 78372 173540 78428
rect 173596 78372 173644 78428
rect 173700 78372 173710 78428
rect 4466 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4750 77644
rect 35186 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35470 77644
rect 65906 77588 65916 77644
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 66180 77588 66190 77644
rect 96626 77588 96636 77644
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96900 77588 96910 77644
rect 127346 77588 127356 77644
rect 127412 77588 127460 77644
rect 127516 77588 127564 77644
rect 127620 77588 127630 77644
rect 158066 77588 158076 77644
rect 158132 77588 158180 77644
rect 158236 77588 158284 77644
rect 158340 77588 158350 77644
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 81266 76804 81276 76860
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81540 76804 81550 76860
rect 111986 76804 111996 76860
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 112260 76804 112270 76860
rect 142706 76804 142716 76860
rect 142772 76804 142820 76860
rect 142876 76804 142924 76860
rect 142980 76804 142990 76860
rect 173426 76804 173436 76860
rect 173492 76804 173540 76860
rect 173596 76804 173644 76860
rect 173700 76804 173710 76860
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 96626 76020 96636 76076
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96900 76020 96910 76076
rect 127346 76020 127356 76076
rect 127412 76020 127460 76076
rect 127516 76020 127564 76076
rect 127620 76020 127630 76076
rect 158066 76020 158076 76076
rect 158132 76020 158180 76076
rect 158236 76020 158284 76076
rect 158340 76020 158350 76076
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 81266 75236 81276 75292
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81540 75236 81550 75292
rect 111986 75236 111996 75292
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 112260 75236 112270 75292
rect 142706 75236 142716 75292
rect 142772 75236 142820 75292
rect 142876 75236 142924 75292
rect 142980 75236 142990 75292
rect 173426 75236 173436 75292
rect 173492 75236 173540 75292
rect 173596 75236 173644 75292
rect 173700 75236 173710 75292
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 96626 74452 96636 74508
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96900 74452 96910 74508
rect 127346 74452 127356 74508
rect 127412 74452 127460 74508
rect 127516 74452 127564 74508
rect 127620 74452 127630 74508
rect 158066 74452 158076 74508
rect 158132 74452 158180 74508
rect 158236 74452 158284 74508
rect 158340 74452 158350 74508
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 81266 73668 81276 73724
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81540 73668 81550 73724
rect 111986 73668 111996 73724
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 112260 73668 112270 73724
rect 142706 73668 142716 73724
rect 142772 73668 142820 73724
rect 142876 73668 142924 73724
rect 142980 73668 142990 73724
rect 173426 73668 173436 73724
rect 173492 73668 173540 73724
rect 173596 73668 173644 73724
rect 173700 73668 173710 73724
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 96626 72884 96636 72940
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96900 72884 96910 72940
rect 127346 72884 127356 72940
rect 127412 72884 127460 72940
rect 127516 72884 127564 72940
rect 127620 72884 127630 72940
rect 158066 72884 158076 72940
rect 158132 72884 158180 72940
rect 158236 72884 158284 72940
rect 158340 72884 158350 72940
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 81266 72100 81276 72156
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81540 72100 81550 72156
rect 111986 72100 111996 72156
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 112260 72100 112270 72156
rect 142706 72100 142716 72156
rect 142772 72100 142820 72156
rect 142876 72100 142924 72156
rect 142980 72100 142990 72156
rect 173426 72100 173436 72156
rect 173492 72100 173540 72156
rect 173596 72100 173644 72156
rect 173700 72100 173710 72156
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 96626 71316 96636 71372
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96900 71316 96910 71372
rect 127346 71316 127356 71372
rect 127412 71316 127460 71372
rect 127516 71316 127564 71372
rect 127620 71316 127630 71372
rect 158066 71316 158076 71372
rect 158132 71316 158180 71372
rect 158236 71316 158284 71372
rect 158340 71316 158350 71372
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 81266 70532 81276 70588
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81540 70532 81550 70588
rect 111986 70532 111996 70588
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 112260 70532 112270 70588
rect 142706 70532 142716 70588
rect 142772 70532 142820 70588
rect 142876 70532 142924 70588
rect 142980 70532 142990 70588
rect 173426 70532 173436 70588
rect 173492 70532 173540 70588
rect 173596 70532 173644 70588
rect 173700 70532 173710 70588
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 96626 69748 96636 69804
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96900 69748 96910 69804
rect 127346 69748 127356 69804
rect 127412 69748 127460 69804
rect 127516 69748 127564 69804
rect 127620 69748 127630 69804
rect 158066 69748 158076 69804
rect 158132 69748 158180 69804
rect 158236 69748 158284 69804
rect 158340 69748 158350 69804
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 81266 68964 81276 69020
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81540 68964 81550 69020
rect 111986 68964 111996 69020
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 112260 68964 112270 69020
rect 142706 68964 142716 69020
rect 142772 68964 142820 69020
rect 142876 68964 142924 69020
rect 142980 68964 142990 69020
rect 173426 68964 173436 69020
rect 173492 68964 173540 69020
rect 173596 68964 173644 69020
rect 173700 68964 173710 69020
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 96626 68180 96636 68236
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96900 68180 96910 68236
rect 127346 68180 127356 68236
rect 127412 68180 127460 68236
rect 127516 68180 127564 68236
rect 127620 68180 127630 68236
rect 158066 68180 158076 68236
rect 158132 68180 158180 68236
rect 158236 68180 158284 68236
rect 158340 68180 158350 68236
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 81266 67396 81276 67452
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81540 67396 81550 67452
rect 111986 67396 111996 67452
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 112260 67396 112270 67452
rect 142706 67396 142716 67452
rect 142772 67396 142820 67452
rect 142876 67396 142924 67452
rect 142980 67396 142990 67452
rect 173426 67396 173436 67452
rect 173492 67396 173540 67452
rect 173596 67396 173644 67452
rect 173700 67396 173710 67452
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 96626 66612 96636 66668
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96900 66612 96910 66668
rect 127346 66612 127356 66668
rect 127412 66612 127460 66668
rect 127516 66612 127564 66668
rect 127620 66612 127630 66668
rect 158066 66612 158076 66668
rect 158132 66612 158180 66668
rect 158236 66612 158284 66668
rect 158340 66612 158350 66668
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 81266 65828 81276 65884
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81540 65828 81550 65884
rect 111986 65828 111996 65884
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 112260 65828 112270 65884
rect 142706 65828 142716 65884
rect 142772 65828 142820 65884
rect 142876 65828 142924 65884
rect 142980 65828 142990 65884
rect 173426 65828 173436 65884
rect 173492 65828 173540 65884
rect 173596 65828 173644 65884
rect 173700 65828 173710 65884
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 96626 65044 96636 65100
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96900 65044 96910 65100
rect 127346 65044 127356 65100
rect 127412 65044 127460 65100
rect 127516 65044 127564 65100
rect 127620 65044 127630 65100
rect 158066 65044 158076 65100
rect 158132 65044 158180 65100
rect 158236 65044 158284 65100
rect 158340 65044 158350 65100
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 81266 64260 81276 64316
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81540 64260 81550 64316
rect 111986 64260 111996 64316
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 112260 64260 112270 64316
rect 142706 64260 142716 64316
rect 142772 64260 142820 64316
rect 142876 64260 142924 64316
rect 142980 64260 142990 64316
rect 173426 64260 173436 64316
rect 173492 64260 173540 64316
rect 173596 64260 173644 64316
rect 173700 64260 173710 64316
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 96626 63476 96636 63532
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96900 63476 96910 63532
rect 127346 63476 127356 63532
rect 127412 63476 127460 63532
rect 127516 63476 127564 63532
rect 127620 63476 127630 63532
rect 158066 63476 158076 63532
rect 158132 63476 158180 63532
rect 158236 63476 158284 63532
rect 158340 63476 158350 63532
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 81266 62692 81276 62748
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81540 62692 81550 62748
rect 111986 62692 111996 62748
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 112260 62692 112270 62748
rect 142706 62692 142716 62748
rect 142772 62692 142820 62748
rect 142876 62692 142924 62748
rect 142980 62692 142990 62748
rect 173426 62692 173436 62748
rect 173492 62692 173540 62748
rect 173596 62692 173644 62748
rect 173700 62692 173710 62748
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 96626 61908 96636 61964
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96900 61908 96910 61964
rect 127346 61908 127356 61964
rect 127412 61908 127460 61964
rect 127516 61908 127564 61964
rect 127620 61908 127630 61964
rect 158066 61908 158076 61964
rect 158132 61908 158180 61964
rect 158236 61908 158284 61964
rect 158340 61908 158350 61964
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 81266 61124 81276 61180
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81540 61124 81550 61180
rect 111986 61124 111996 61180
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 112260 61124 112270 61180
rect 142706 61124 142716 61180
rect 142772 61124 142820 61180
rect 142876 61124 142924 61180
rect 142980 61124 142990 61180
rect 173426 61124 173436 61180
rect 173492 61124 173540 61180
rect 173596 61124 173644 61180
rect 173700 61124 173710 61180
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 96626 60340 96636 60396
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96900 60340 96910 60396
rect 127346 60340 127356 60396
rect 127412 60340 127460 60396
rect 127516 60340 127564 60396
rect 127620 60340 127630 60396
rect 158066 60340 158076 60396
rect 158132 60340 158180 60396
rect 158236 60340 158284 60396
rect 158340 60340 158350 60396
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 81266 59556 81276 59612
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81540 59556 81550 59612
rect 111986 59556 111996 59612
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 112260 59556 112270 59612
rect 142706 59556 142716 59612
rect 142772 59556 142820 59612
rect 142876 59556 142924 59612
rect 142980 59556 142990 59612
rect 173426 59556 173436 59612
rect 173492 59556 173540 59612
rect 173596 59556 173644 59612
rect 173700 59556 173710 59612
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 96626 58772 96636 58828
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96900 58772 96910 58828
rect 127346 58772 127356 58828
rect 127412 58772 127460 58828
rect 127516 58772 127564 58828
rect 127620 58772 127630 58828
rect 158066 58772 158076 58828
rect 158132 58772 158180 58828
rect 158236 58772 158284 58828
rect 158340 58772 158350 58828
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 81266 57988 81276 58044
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81540 57988 81550 58044
rect 111986 57988 111996 58044
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 112260 57988 112270 58044
rect 142706 57988 142716 58044
rect 142772 57988 142820 58044
rect 142876 57988 142924 58044
rect 142980 57988 142990 58044
rect 173426 57988 173436 58044
rect 173492 57988 173540 58044
rect 173596 57988 173644 58044
rect 173700 57988 173710 58044
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 96626 57204 96636 57260
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96900 57204 96910 57260
rect 127346 57204 127356 57260
rect 127412 57204 127460 57260
rect 127516 57204 127564 57260
rect 127620 57204 127630 57260
rect 158066 57204 158076 57260
rect 158132 57204 158180 57260
rect 158236 57204 158284 57260
rect 158340 57204 158350 57260
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 81266 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81550 56476
rect 111986 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112270 56476
rect 142706 56420 142716 56476
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142980 56420 142990 56476
rect 173426 56420 173436 56476
rect 173492 56420 173540 56476
rect 173596 56420 173644 56476
rect 173700 56420 173710 56476
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 96626 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96910 55692
rect 127346 55636 127356 55692
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127620 55636 127630 55692
rect 158066 55636 158076 55692
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158340 55636 158350 55692
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 81266 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81550 54908
rect 111986 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112270 54908
rect 142706 54852 142716 54908
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142980 54852 142990 54908
rect 173426 54852 173436 54908
rect 173492 54852 173540 54908
rect 173596 54852 173644 54908
rect 173700 54852 173710 54908
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 96626 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96910 54124
rect 127346 54068 127356 54124
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127620 54068 127630 54124
rect 158066 54068 158076 54124
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158340 54068 158350 54124
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 81266 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81550 53340
rect 111986 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112270 53340
rect 142706 53284 142716 53340
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142980 53284 142990 53340
rect 173426 53284 173436 53340
rect 173492 53284 173540 53340
rect 173596 53284 173644 53340
rect 173700 53284 173710 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 96626 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96910 52556
rect 127346 52500 127356 52556
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127620 52500 127630 52556
rect 158066 52500 158076 52556
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158340 52500 158350 52556
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 81266 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81550 51772
rect 111986 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112270 51772
rect 142706 51716 142716 51772
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142980 51716 142990 51772
rect 173426 51716 173436 51772
rect 173492 51716 173540 51772
rect 173596 51716 173644 51772
rect 173700 51716 173710 51772
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 96626 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96910 50988
rect 127346 50932 127356 50988
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127620 50932 127630 50988
rect 158066 50932 158076 50988
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158340 50932 158350 50988
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 81266 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81550 50204
rect 111986 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112270 50204
rect 142706 50148 142716 50204
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142980 50148 142990 50204
rect 173426 50148 173436 50204
rect 173492 50148 173540 50204
rect 173596 50148 173644 50204
rect 173700 50148 173710 50204
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 96626 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96910 49420
rect 127346 49364 127356 49420
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127620 49364 127630 49420
rect 158066 49364 158076 49420
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158340 49364 158350 49420
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 81266 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81550 48636
rect 111986 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112270 48636
rect 142706 48580 142716 48636
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142980 48580 142990 48636
rect 173426 48580 173436 48636
rect 173492 48580 173540 48636
rect 173596 48580 173644 48636
rect 173700 48580 173710 48636
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 96626 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96910 47852
rect 127346 47796 127356 47852
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127620 47796 127630 47852
rect 158066 47796 158076 47852
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158340 47796 158350 47852
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 81266 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81550 47068
rect 111986 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112270 47068
rect 142706 47012 142716 47068
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142980 47012 142990 47068
rect 173426 47012 173436 47068
rect 173492 47012 173540 47068
rect 173596 47012 173644 47068
rect 173700 47012 173710 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 96626 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96910 46284
rect 127346 46228 127356 46284
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127620 46228 127630 46284
rect 158066 46228 158076 46284
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158340 46228 158350 46284
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 81266 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81550 45500
rect 111986 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112270 45500
rect 142706 45444 142716 45500
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142980 45444 142990 45500
rect 173426 45444 173436 45500
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173700 45444 173710 45500
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 96626 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96910 44716
rect 127346 44660 127356 44716
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127620 44660 127630 44716
rect 158066 44660 158076 44716
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158340 44660 158350 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 81266 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81550 43932
rect 111986 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112270 43932
rect 142706 43876 142716 43932
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142980 43876 142990 43932
rect 173426 43876 173436 43932
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173700 43876 173710 43932
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 96626 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96910 43148
rect 127346 43092 127356 43148
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127620 43092 127630 43148
rect 158066 43092 158076 43148
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158340 43092 158350 43148
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 81266 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81550 42364
rect 111986 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112270 42364
rect 142706 42308 142716 42364
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142980 42308 142990 42364
rect 173426 42308 173436 42364
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173700 42308 173710 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 96626 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96910 41580
rect 127346 41524 127356 41580
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127620 41524 127630 41580
rect 158066 41524 158076 41580
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158340 41524 158350 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 81266 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81550 40796
rect 111986 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112270 40796
rect 142706 40740 142716 40796
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142980 40740 142990 40796
rect 173426 40740 173436 40796
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173700 40740 173710 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 96626 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96910 40012
rect 127346 39956 127356 40012
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127620 39956 127630 40012
rect 158066 39956 158076 40012
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158340 39956 158350 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 81266 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81550 39228
rect 111986 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112270 39228
rect 142706 39172 142716 39228
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142980 39172 142990 39228
rect 173426 39172 173436 39228
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173700 39172 173710 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 96626 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96910 38444
rect 127346 38388 127356 38444
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127620 38388 127630 38444
rect 158066 38388 158076 38444
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158340 38388 158350 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 81266 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81550 37660
rect 111986 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112270 37660
rect 142706 37604 142716 37660
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142980 37604 142990 37660
rect 173426 37604 173436 37660
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173700 37604 173710 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 96626 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96910 36876
rect 127346 36820 127356 36876
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127620 36820 127630 36876
rect 158066 36820 158076 36876
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158340 36820 158350 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 81266 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81550 36092
rect 111986 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112270 36092
rect 142706 36036 142716 36092
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142980 36036 142990 36092
rect 173426 36036 173436 36092
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173700 36036 173710 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 96626 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96910 35308
rect 127346 35252 127356 35308
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127620 35252 127630 35308
rect 158066 35252 158076 35308
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158340 35252 158350 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 81266 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81550 34524
rect 111986 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112270 34524
rect 142706 34468 142716 34524
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142980 34468 142990 34524
rect 173426 34468 173436 34524
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173700 34468 173710 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 96626 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96910 33740
rect 127346 33684 127356 33740
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127620 33684 127630 33740
rect 158066 33684 158076 33740
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158340 33684 158350 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 81266 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81550 32956
rect 111986 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112270 32956
rect 142706 32900 142716 32956
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142980 32900 142990 32956
rect 173426 32900 173436 32956
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173700 32900 173710 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 96626 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96910 32172
rect 127346 32116 127356 32172
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127620 32116 127630 32172
rect 158066 32116 158076 32172
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158340 32116 158350 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 81266 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81550 31388
rect 111986 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112270 31388
rect 142706 31332 142716 31388
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142980 31332 142990 31388
rect 173426 31332 173436 31388
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173700 31332 173710 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 96626 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96910 30604
rect 127346 30548 127356 30604
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127620 30548 127630 30604
rect 158066 30548 158076 30604
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158340 30548 158350 30604
rect 49186 30268 49196 30324
rect 49252 30268 102396 30324
rect 102452 30268 102462 30324
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 81266 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81550 29820
rect 111986 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112270 29820
rect 142706 29764 142716 29820
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142980 29764 142990 29820
rect 173426 29764 173436 29820
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173700 29764 173710 29820
rect 43698 29372 43708 29428
rect 43764 29372 74844 29428
rect 74900 29372 74910 29428
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 96626 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96910 29036
rect 127346 28980 127356 29036
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127620 28980 127630 29036
rect 158066 28980 158076 29036
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158340 28980 158350 29036
rect 70130 28588 70140 28644
rect 70196 28588 126364 28644
rect 126420 28588 126430 28644
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 81266 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81550 28252
rect 111986 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112270 28252
rect 142706 28196 142716 28252
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142980 28196 142990 28252
rect 173426 28196 173436 28252
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173700 28196 173710 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 96626 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96910 27468
rect 127346 27412 127356 27468
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127620 27412 127630 27468
rect 158066 27412 158076 27468
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158340 27412 158350 27468
rect 67890 27356 67900 27412
rect 67956 27356 71372 27412
rect 71428 27356 71438 27412
rect 45266 27244 45276 27300
rect 45332 27244 97468 27300
rect 97524 27244 98364 27300
rect 98420 27244 98430 27300
rect 45714 27132 45724 27188
rect 45780 27132 108668 27188
rect 108724 27132 108734 27188
rect 41010 27020 41020 27076
rect 41076 27020 120540 27076
rect 120596 27020 120606 27076
rect 40002 26908 40012 26964
rect 40068 26908 120764 26964
rect 120820 26908 120830 26964
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 81266 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81550 26684
rect 111986 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112270 26684
rect 142706 26628 142716 26684
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142980 26628 142990 26684
rect 173426 26628 173436 26684
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173700 26628 173710 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 96626 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96910 25900
rect 127346 25844 127356 25900
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127620 25844 127630 25900
rect 158066 25844 158076 25900
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158340 25844 158350 25900
rect 40226 25564 40236 25620
rect 40292 25564 90860 25620
rect 90916 25564 91532 25620
rect 91588 25564 91598 25620
rect 52770 25452 52780 25508
rect 52836 25452 104412 25508
rect 104468 25452 104478 25508
rect 68786 25340 68796 25396
rect 68852 25340 124236 25396
rect 124292 25340 124302 25396
rect 72146 25228 72156 25284
rect 72212 25228 127708 25284
rect 127764 25228 127774 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 81266 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81550 25116
rect 111986 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112270 25116
rect 142706 25060 142716 25116
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142980 25060 142990 25116
rect 173426 25060 173436 25116
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173700 25060 173710 25116
rect 100706 24444 100716 24500
rect 100772 24444 169148 24500
rect 169204 24444 169214 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 96626 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96910 24332
rect 127346 24276 127356 24332
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127620 24276 127630 24332
rect 158066 24276 158076 24332
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158340 24276 158350 24332
rect 65538 24108 65548 24164
rect 65604 24108 118300 24164
rect 118356 24108 118366 24164
rect 70242 23996 70252 24052
rect 70308 23996 124572 24052
rect 124628 23996 124638 24052
rect 78866 23884 78876 23940
rect 78932 23884 133980 23940
rect 134036 23884 134046 23940
rect 48626 23772 48636 23828
rect 48692 23772 106092 23828
rect 106148 23772 106158 23828
rect 46946 23660 46956 23716
rect 47012 23660 112364 23716
rect 112420 23660 112430 23716
rect 52882 23548 52892 23604
rect 52948 23548 53564 23604
rect 53620 23548 79436 23604
rect 79492 23548 79502 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 81266 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81550 23548
rect 111986 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112270 23548
rect 142706 23492 142716 23548
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142980 23492 142990 23548
rect 173426 23492 173436 23548
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173700 23492 173710 23548
rect 38546 22988 38556 23044
rect 38612 22988 80780 23044
rect 80836 22988 81116 23044
rect 81172 22988 81182 23044
rect 44706 22876 44716 22932
rect 44772 22876 113148 22932
rect 113204 22876 113214 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 96626 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96910 22764
rect 127346 22708 127356 22764
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127620 22708 127630 22764
rect 158066 22708 158076 22764
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158340 22708 158350 22764
rect 69906 22652 69916 22708
rect 69972 22652 83916 22708
rect 83972 22652 83982 22708
rect 25778 22540 25788 22596
rect 25844 22540 84476 22596
rect 84532 22540 84542 22596
rect 33618 22428 33628 22484
rect 33684 22428 34860 22484
rect 34916 22428 43708 22484
rect 74722 22428 74732 22484
rect 74788 22428 135548 22484
rect 135604 22428 135614 22484
rect 43652 22260 43708 22428
rect 74946 22316 74956 22372
rect 75012 22316 133532 22372
rect 133588 22316 133598 22372
rect 43652 22204 73948 22260
rect 74004 22204 74014 22260
rect 82002 22204 82012 22260
rect 82068 22204 123340 22260
rect 123396 22204 123406 22260
rect 69682 22092 69692 22148
rect 69748 22092 130396 22148
rect 130452 22092 130462 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 81266 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81550 21980
rect 111986 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112270 21980
rect 142706 21924 142716 21980
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142980 21924 142990 21980
rect 173426 21924 173436 21980
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173700 21924 173710 21980
rect 58146 21420 58156 21476
rect 58212 21420 102060 21476
rect 102116 21420 102126 21476
rect 46274 21308 46284 21364
rect 46340 21308 104300 21364
rect 104356 21308 104366 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 96626 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96910 21196
rect 127346 21140 127356 21196
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127620 21140 127630 21196
rect 158066 21140 158076 21196
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158340 21140 158350 21196
rect 48738 20972 48748 21028
rect 48804 20972 76076 21028
rect 76132 20972 76142 21028
rect 99026 20860 99036 20916
rect 99092 20860 167356 20916
rect 167412 20860 167422 20916
rect 77858 20748 77868 20804
rect 77924 20748 115052 20804
rect 115108 20748 115118 20804
rect 84802 20636 84812 20692
rect 84868 20636 127148 20692
rect 127204 20636 127214 20692
rect 71250 20524 71260 20580
rect 71316 20524 123676 20580
rect 123732 20524 123742 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 81266 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81550 20412
rect 111986 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112270 20412
rect 142706 20356 142716 20412
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142980 20356 142990 20412
rect 173426 20356 173436 20412
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173700 20356 173710 20412
rect 8978 20188 8988 20244
rect 9044 20188 128492 20244
rect 128548 20188 128558 20244
rect 68226 19740 68236 19796
rect 68292 19740 114828 19796
rect 114884 19740 114894 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 96626 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96910 19628
rect 127346 19572 127356 19628
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127620 19572 127630 19628
rect 158066 19572 158076 19628
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158340 19572 158350 19628
rect 35074 19404 35084 19460
rect 35140 19404 62860 19460
rect 62916 19404 81004 19460
rect 81060 19404 81070 19460
rect 12562 19292 12572 19348
rect 12628 19292 63756 19348
rect 63812 19292 63822 19348
rect 66994 19292 67004 19348
rect 67060 19292 113596 19348
rect 113652 19292 113662 19348
rect 115826 19292 115836 19348
rect 115892 19292 140700 19348
rect 140756 19292 140766 19348
rect 86930 19180 86940 19236
rect 86996 19180 125692 19236
rect 125748 19180 125758 19236
rect 57026 19068 57036 19124
rect 57092 19068 94444 19124
rect 94500 19068 94510 19124
rect 95554 19068 95564 19124
rect 95620 19068 135772 19124
rect 135828 19068 135838 19124
rect 58482 18956 58492 19012
rect 58548 18956 101276 19012
rect 101332 18956 101342 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 81266 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81550 18844
rect 111986 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112270 18844
rect 142706 18788 142716 18844
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142980 18788 142990 18844
rect 173426 18788 173436 18844
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173700 18788 173710 18844
rect 23090 18620 23100 18676
rect 23156 18620 82348 18676
rect 82404 18620 82414 18676
rect 85922 18620 85932 18676
rect 85988 18620 134764 18676
rect 134820 18620 134830 18676
rect 16818 18508 16828 18564
rect 16884 18508 78204 18564
rect 78260 18508 78270 18564
rect 107090 18508 107100 18564
rect 107156 18508 163436 18564
rect 163492 18508 163502 18564
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 96626 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96910 18060
rect 127346 18004 127356 18060
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127620 18004 127630 18060
rect 158066 18004 158076 18060
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158340 18004 158350 18060
rect 92194 17836 92204 17892
rect 92260 17836 137228 17892
rect 137284 17836 137294 17892
rect 87042 17724 87052 17780
rect 87108 17724 136780 17780
rect 136836 17724 136846 17780
rect 32946 17612 32956 17668
rect 33012 17612 88844 17668
rect 88900 17612 88910 17668
rect 114146 17612 114156 17668
rect 114212 17612 136892 17668
rect 136948 17612 136958 17668
rect 46834 17500 46844 17556
rect 46900 17500 123228 17556
rect 123284 17500 123294 17556
rect 62178 17388 62188 17444
rect 62244 17388 95676 17444
rect 95732 17388 95742 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 81266 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81550 17276
rect 111986 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112270 17276
rect 142706 17220 142716 17276
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142980 17220 142990 17276
rect 173426 17220 173436 17276
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173700 17220 173710 17276
rect 47954 17052 47964 17108
rect 48020 17052 114268 17108
rect 114324 17052 114334 17108
rect 48962 16940 48972 16996
rect 49028 16940 121212 16996
rect 121268 16940 121278 16996
rect 15138 16828 15148 16884
rect 15204 16828 80556 16884
rect 80612 16828 80622 16884
rect 97570 16828 97580 16884
rect 97636 16828 113260 16884
rect 113316 16828 114268 16884
rect 114212 16772 114268 16828
rect 26898 16716 26908 16772
rect 26964 16716 33628 16772
rect 33684 16716 33694 16772
rect 114212 16716 131740 16772
rect 131796 16716 131806 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 96626 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96910 16492
rect 127346 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127630 16492
rect 158066 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158350 16492
rect 63410 16268 63420 16324
rect 63476 16268 95228 16324
rect 95284 16268 95294 16324
rect 58930 16156 58940 16212
rect 58996 16156 94780 16212
rect 94836 16156 94846 16212
rect 29698 16044 29708 16100
rect 29764 16044 89852 16100
rect 89908 16044 89918 16100
rect 57698 15932 57708 15988
rect 57764 15932 96348 15988
rect 96404 15932 96414 15988
rect 43026 15820 43036 15876
rect 43092 15820 77644 15876
rect 77700 15820 77710 15876
rect 97122 15820 97132 15876
rect 97188 15820 116396 15876
rect 116452 15820 116462 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 81266 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81550 15708
rect 111986 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112270 15708
rect 142706 15652 142716 15708
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142980 15652 142990 15708
rect 173426 15652 173436 15708
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173700 15652 173710 15708
rect 93426 15484 93436 15540
rect 93492 15484 131516 15540
rect 131572 15484 131582 15540
rect 37874 15372 37884 15428
rect 37940 15372 87836 15428
rect 87892 15372 87902 15428
rect 92306 15372 92316 15428
rect 92372 15372 142604 15428
rect 142660 15372 142670 15428
rect 72930 15260 72940 15316
rect 72996 15260 128156 15316
rect 128212 15260 128222 15316
rect 85586 15148 85596 15204
rect 85652 15148 137004 15204
rect 137060 15148 137070 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 96626 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96910 14924
rect 127346 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127630 14924
rect 158066 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158350 14924
rect 61730 14700 61740 14756
rect 61796 14700 93996 14756
rect 94052 14700 94062 14756
rect 55794 14588 55804 14644
rect 55860 14588 105756 14644
rect 105812 14588 105822 14644
rect 60498 14476 60508 14532
rect 60564 14476 100604 14532
rect 100660 14476 100670 14532
rect 74050 14364 74060 14420
rect 74116 14364 115276 14420
rect 115332 14364 115342 14420
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 81266 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81550 14140
rect 111986 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112270 14140
rect 142706 14084 142716 14140
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142980 14084 142990 14140
rect 173426 14084 173436 14140
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173700 14084 173710 14140
rect 106866 14028 106876 14084
rect 106932 14028 111804 14084
rect 111860 14028 111870 14084
rect 56578 13916 56588 13972
rect 56644 13916 94108 13972
rect 94164 13916 94174 13972
rect 100482 13916 100492 13972
rect 100548 13916 137116 13972
rect 137172 13916 137182 13972
rect 77298 13804 77308 13860
rect 77364 13804 85708 13860
rect 91746 13804 91756 13860
rect 91812 13804 141820 13860
rect 141876 13804 141886 13860
rect 28466 13692 28476 13748
rect 28532 13692 79884 13748
rect 79940 13692 79950 13748
rect 21970 13580 21980 13636
rect 22036 13580 61516 13636
rect 61572 13580 61582 13636
rect 68338 13580 68348 13636
rect 68404 13580 68796 13636
rect 68852 13580 69132 13636
rect 69188 13580 69198 13636
rect 69570 13580 69580 13636
rect 69636 13580 71372 13636
rect 71428 13580 72716 13636
rect 72772 13580 72782 13636
rect 77074 13580 77084 13636
rect 77140 13580 77420 13636
rect 77476 13580 77486 13636
rect 78642 13580 78652 13636
rect 78708 13580 78876 13636
rect 78932 13580 79100 13636
rect 79156 13580 79166 13636
rect 85652 13524 85708 13804
rect 91522 13692 91532 13748
rect 91588 13692 141372 13748
rect 141428 13692 141438 13748
rect 109218 13580 109228 13636
rect 109284 13580 111580 13636
rect 111636 13580 111646 13636
rect 111794 13580 111804 13636
rect 111860 13580 161308 13636
rect 161364 13580 161374 13636
rect 73938 13468 73948 13524
rect 74004 13468 75404 13524
rect 75460 13468 75628 13524
rect 75684 13468 75694 13524
rect 77186 13468 77196 13524
rect 77252 13468 78764 13524
rect 78820 13468 78830 13524
rect 80210 13468 80220 13524
rect 80276 13468 83020 13524
rect 83076 13468 83086 13524
rect 85652 13468 133756 13524
rect 133812 13468 133822 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 96626 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96910 13356
rect 127346 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127630 13356
rect 158066 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158350 13356
rect 55412 13132 77084 13188
rect 77140 13132 77150 13188
rect 55412 12852 55468 13132
rect 69346 13020 69356 13076
rect 69412 13020 70140 13076
rect 70196 13020 70206 13076
rect 74834 13020 74844 13076
rect 74900 13020 76524 13076
rect 76580 13020 77420 13076
rect 77476 13020 77486 13076
rect 83010 13020 83020 13076
rect 83076 13020 85372 13076
rect 85428 13020 85438 13076
rect 71026 12908 71036 12964
rect 71092 12908 71484 12964
rect 71540 12908 71550 12964
rect 76626 12908 76636 12964
rect 76692 12908 79716 12964
rect 82114 12908 82124 12964
rect 82180 12908 143724 12964
rect 143780 12908 143790 12964
rect 79660 12852 79716 12908
rect 24434 12796 24444 12852
rect 24500 12796 55468 12852
rect 68450 12796 68460 12852
rect 68516 12796 75964 12852
rect 76020 12796 77084 12852
rect 77140 12796 77150 12852
rect 79650 12796 79660 12852
rect 79716 12796 79884 12852
rect 79940 12796 82012 12852
rect 82068 12796 82078 12852
rect 74722 12684 74732 12740
rect 74788 12684 75180 12740
rect 75236 12684 75246 12740
rect 79426 12684 79436 12740
rect 79492 12684 81116 12740
rect 81172 12684 81452 12740
rect 81508 12684 81518 12740
rect 100370 12684 100380 12740
rect 100436 12684 101164 12740
rect 101220 12684 101230 12740
rect 107202 12684 107212 12740
rect 107268 12684 129836 12740
rect 129892 12684 129902 12740
rect 55412 12572 76188 12628
rect 76244 12572 76254 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 55412 12516 55468 12572
rect 81266 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81550 12572
rect 111986 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112270 12572
rect 142706 12516 142716 12572
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142980 12516 142990 12572
rect 173426 12516 173436 12572
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173700 12516 173710 12572
rect 51538 12460 51548 12516
rect 51604 12460 55468 12516
rect 56242 12460 56252 12516
rect 56308 12460 57036 12516
rect 57092 12460 57932 12516
rect 57988 12460 57998 12516
rect 70914 12460 70924 12516
rect 70980 12460 72156 12516
rect 72212 12460 72222 12516
rect 74946 12460 74956 12516
rect 75012 12460 78540 12516
rect 78596 12460 79996 12516
rect 80052 12460 80556 12516
rect 80612 12460 80622 12516
rect 80556 12404 80612 12460
rect 36866 12348 36876 12404
rect 36932 12348 68460 12404
rect 68516 12348 68526 12404
rect 70214 12348 70252 12404
rect 70308 12348 70318 12404
rect 72258 12348 72268 12404
rect 72324 12348 74172 12404
rect 74228 12348 74238 12404
rect 75842 12348 75852 12404
rect 75908 12348 76076 12404
rect 76132 12348 76142 12404
rect 77074 12348 77084 12404
rect 77140 12348 77980 12404
rect 78036 12348 78046 12404
rect 80556 12348 81676 12404
rect 81732 12348 81742 12404
rect 82002 12348 82012 12404
rect 82068 12348 82572 12404
rect 82628 12348 82638 12404
rect 114706 12348 114716 12404
rect 114772 12348 142492 12404
rect 142548 12348 142558 12404
rect 57362 12236 57372 12292
rect 57428 12236 58604 12292
rect 58660 12236 59612 12292
rect 59668 12236 60844 12292
rect 60900 12236 60910 12292
rect 63746 12236 63756 12292
rect 63812 12236 64540 12292
rect 64596 12236 73612 12292
rect 73668 12236 73678 12292
rect 77186 12236 77196 12292
rect 77252 12236 85708 12292
rect 92082 12236 92092 12292
rect 92148 12236 136668 12292
rect 136724 12236 136734 12292
rect 85652 12180 85708 12236
rect 29922 12124 29932 12180
rect 29988 12124 76020 12180
rect 76178 12124 76188 12180
rect 76244 12124 79212 12180
rect 79268 12124 79278 12180
rect 85652 12124 89516 12180
rect 89572 12124 89582 12180
rect 93650 12124 93660 12180
rect 93716 12124 145964 12180
rect 146020 12124 146030 12180
rect 75964 12068 76020 12124
rect 59154 12012 59164 12068
rect 59220 12012 61180 12068
rect 61236 12012 61246 12068
rect 65426 12012 65436 12068
rect 65492 12012 66108 12068
rect 66164 12012 66892 12068
rect 66948 12012 66958 12068
rect 69794 12012 69804 12068
rect 69860 12012 70028 12068
rect 70084 12012 70588 12068
rect 70644 12012 71036 12068
rect 71092 12012 71102 12068
rect 73042 12012 73052 12068
rect 73108 12012 75740 12068
rect 75796 12012 75806 12068
rect 75964 12012 76972 12068
rect 77028 12012 77038 12068
rect 77410 12012 77420 12068
rect 77476 12012 80108 12068
rect 80164 12012 80174 12068
rect 82226 12012 82236 12068
rect 82292 12012 83356 12068
rect 83412 12012 83422 12068
rect 105410 12012 105420 12068
rect 105476 12012 105980 12068
rect 106036 12012 106046 12068
rect 106754 12012 106764 12068
rect 106820 12012 108108 12068
rect 108164 12012 108174 12068
rect 109442 12012 109452 12068
rect 109508 12012 112140 12068
rect 112196 12012 117180 12068
rect 117236 12012 117246 12068
rect 129266 12012 129276 12068
rect 129332 12012 161420 12068
rect 161476 12012 161486 12068
rect 60610 11900 60620 11956
rect 60676 11900 61964 11956
rect 62020 11900 90188 11956
rect 90244 11900 90254 11956
rect 100258 11900 100268 11956
rect 100324 11900 104076 11956
rect 104132 11900 110628 11956
rect 51986 11788 51996 11844
rect 52052 11788 52892 11844
rect 52948 11788 52958 11844
rect 71026 11788 71036 11844
rect 71092 11788 74508 11844
rect 74564 11788 74574 11844
rect 78306 11788 78316 11844
rect 78372 11788 79100 11844
rect 79156 11788 79660 11844
rect 79716 11788 80892 11844
rect 80948 11788 80958 11844
rect 81330 11788 81340 11844
rect 81396 11788 82348 11844
rect 82404 11788 83244 11844
rect 83300 11788 83310 11844
rect 91522 11788 91532 11844
rect 91588 11788 93548 11844
rect 93604 11788 93614 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 96626 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96910 11788
rect 110572 11732 110628 11900
rect 111244 11900 170380 11956
rect 170436 11900 170446 11956
rect 111244 11844 111300 11900
rect 110786 11788 110796 11844
rect 110852 11788 111300 11844
rect 111570 11788 111580 11844
rect 111636 11788 112588 11844
rect 112644 11788 112654 11844
rect 115490 11788 115500 11844
rect 115556 11788 120092 11844
rect 120148 11788 120158 11844
rect 115500 11732 115556 11788
rect 127346 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127630 11788
rect 158066 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158350 11788
rect 69122 11676 69132 11732
rect 69188 11676 69692 11732
rect 69748 11676 69758 11732
rect 71586 11676 71596 11732
rect 71652 11676 71932 11732
rect 71988 11676 71998 11732
rect 90402 11676 90412 11732
rect 90468 11676 91084 11732
rect 91140 11676 91150 11732
rect 97122 11676 97132 11732
rect 97188 11676 97692 11732
rect 97748 11676 97758 11732
rect 98130 11676 98140 11732
rect 98196 11676 98812 11732
rect 98868 11676 100156 11732
rect 100212 11676 100222 11732
rect 110572 11676 115556 11732
rect 46162 11564 46172 11620
rect 46228 11564 46956 11620
rect 47012 11564 47022 11620
rect 56130 11564 56140 11620
rect 56196 11564 97020 11620
rect 97076 11564 97086 11620
rect 59378 11452 59388 11508
rect 59444 11452 59948 11508
rect 60004 11452 60508 11508
rect 60564 11452 60574 11508
rect 63718 11452 63756 11508
rect 63812 11452 63822 11508
rect 70130 11452 70140 11508
rect 70196 11452 70812 11508
rect 70868 11452 70878 11508
rect 74162 11452 74172 11508
rect 74228 11452 77196 11508
rect 77252 11452 77262 11508
rect 77522 11452 77532 11508
rect 77588 11452 78092 11508
rect 78148 11452 78158 11508
rect 78530 11452 78540 11508
rect 78596 11452 79324 11508
rect 79380 11452 79390 11508
rect 82114 11452 82124 11508
rect 82180 11452 82796 11508
rect 82852 11452 83468 11508
rect 83524 11452 90412 11508
rect 90468 11452 90478 11508
rect 104290 11452 104300 11508
rect 104356 11452 104748 11508
rect 104804 11452 104814 11508
rect 109172 11452 128044 11508
rect 128100 11452 128110 11508
rect 109172 11396 109228 11452
rect 43250 11340 43260 11396
rect 43316 11340 63980 11396
rect 64036 11340 64046 11396
rect 68562 11340 68572 11396
rect 68628 11340 69692 11396
rect 69748 11340 70028 11396
rect 70084 11340 70700 11396
rect 70756 11340 71708 11396
rect 71764 11340 71774 11396
rect 75730 11340 75740 11396
rect 75796 11340 78204 11396
rect 78260 11340 78428 11396
rect 78484 11340 78494 11396
rect 88946 11340 88956 11396
rect 89012 11340 92428 11396
rect 92484 11340 93772 11396
rect 93828 11340 94220 11396
rect 94276 11340 96460 11396
rect 96516 11340 98140 11396
rect 98196 11340 98206 11396
rect 98924 11340 101052 11396
rect 101108 11340 101118 11396
rect 101714 11340 101724 11396
rect 101780 11340 109228 11396
rect 98924 11284 98980 11340
rect 51090 11228 51100 11284
rect 51156 11228 51324 11284
rect 51380 11228 98980 11284
rect 99148 11228 99932 11284
rect 99988 11228 102508 11284
rect 102564 11228 102574 11284
rect 99148 11172 99204 11228
rect 43138 11116 43148 11172
rect 43204 11116 46620 11172
rect 46676 11116 46686 11172
rect 51650 11116 51660 11172
rect 51716 11116 52780 11172
rect 52836 11116 52846 11172
rect 55458 11116 55468 11172
rect 55524 11116 56028 11172
rect 56084 11116 63196 11172
rect 63252 11116 63262 11172
rect 66546 11116 66556 11172
rect 66612 11116 67116 11172
rect 67172 11116 68124 11172
rect 68180 11116 68572 11172
rect 68628 11116 69244 11172
rect 69300 11116 69310 11172
rect 71586 11116 71596 11172
rect 71652 11116 73276 11172
rect 73332 11116 73342 11172
rect 73490 11116 73500 11172
rect 73556 11116 84476 11172
rect 84532 11116 88396 11172
rect 88452 11116 88462 11172
rect 96002 11116 96012 11172
rect 96068 11116 99148 11172
rect 99204 11116 99214 11172
rect 99810 11116 99820 11172
rect 99876 11116 100716 11172
rect 100772 11116 101164 11172
rect 101220 11116 101230 11172
rect 109890 11116 109900 11172
rect 109956 11116 112756 11172
rect 113138 11116 113148 11172
rect 113204 11116 113260 11172
rect 113316 11116 113326 11172
rect 114678 11116 114716 11172
rect 114772 11116 114782 11172
rect 115266 11116 115276 11172
rect 115332 11116 116732 11172
rect 116788 11116 116798 11172
rect 119298 11116 119308 11172
rect 119364 11116 150444 11172
rect 150500 11116 150510 11172
rect 71596 11060 71652 11116
rect 112700 11060 112756 11116
rect 62626 11004 62636 11060
rect 62692 11004 65660 11060
rect 65716 11004 66332 11060
rect 66388 11004 66398 11060
rect 67442 11004 67452 11060
rect 67508 11004 68684 11060
rect 68740 11004 71652 11060
rect 76178 11004 76188 11060
rect 76244 11004 78316 11060
rect 78372 11004 78382 11060
rect 99474 11004 99484 11060
rect 99540 11004 100044 11060
rect 100100 11004 101500 11060
rect 101556 11004 101566 11060
rect 112690 11004 112700 11060
rect 112756 11004 119084 11060
rect 119140 11004 119150 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 81266 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81550 11004
rect 111986 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112270 11004
rect 142706 10948 142716 11004
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142980 10948 142990 11004
rect 173426 10948 173436 11004
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173700 10948 173710 11004
rect 55412 10892 68572 10948
rect 68628 10892 68638 10948
rect 70130 10892 70140 10948
rect 70196 10892 71260 10948
rect 71316 10892 71326 10948
rect 86370 10892 86380 10948
rect 86436 10892 87612 10948
rect 87668 10892 87678 10948
rect 98242 10892 98252 10948
rect 98308 10892 99036 10948
rect 99092 10892 100380 10948
rect 100436 10892 100446 10948
rect 38546 10780 38556 10836
rect 38612 10780 39340 10836
rect 39396 10780 39406 10836
rect 44930 10780 44940 10836
rect 44996 10780 45276 10836
rect 45332 10780 46396 10836
rect 46452 10780 46462 10836
rect 46610 10780 46620 10836
rect 46676 10780 51100 10836
rect 51156 10780 51166 10836
rect 55412 10724 55468 10892
rect 61506 10780 61516 10836
rect 61572 10780 70252 10836
rect 70308 10780 70318 10836
rect 71148 10780 71484 10836
rect 71540 10780 71550 10836
rect 73826 10780 73836 10836
rect 73892 10780 103628 10836
rect 103684 10780 103694 10836
rect 105746 10780 105756 10836
rect 105812 10780 106428 10836
rect 106484 10780 106494 10836
rect 110450 10780 110460 10836
rect 110516 10780 115892 10836
rect 117394 10780 117404 10836
rect 117460 10780 160412 10836
rect 160468 10780 160478 10836
rect 45042 10668 45052 10724
rect 45108 10668 55468 10724
rect 56914 10668 56924 10724
rect 56980 10668 57484 10724
rect 57540 10668 57550 10724
rect 64866 10668 64876 10724
rect 64932 10668 65996 10724
rect 66052 10668 67340 10724
rect 67396 10668 67406 10724
rect 45714 10556 45724 10612
rect 45780 10556 46620 10612
rect 46676 10556 46686 10612
rect 50866 10556 50876 10612
rect 50932 10556 51884 10612
rect 51940 10556 52668 10612
rect 52724 10556 55916 10612
rect 55972 10556 56812 10612
rect 56868 10556 56878 10612
rect 60498 10556 60508 10612
rect 60564 10556 61628 10612
rect 61684 10556 61694 10612
rect 63970 10556 63980 10612
rect 64036 10556 69244 10612
rect 69300 10556 69310 10612
rect 40898 10444 40908 10500
rect 40964 10444 41580 10500
rect 41636 10444 42700 10500
rect 42756 10444 46060 10500
rect 46116 10444 46732 10500
rect 46788 10444 49868 10500
rect 49924 10444 53564 10500
rect 53620 10444 56140 10500
rect 56196 10444 56476 10500
rect 56532 10444 56542 10500
rect 61180 10444 64764 10500
rect 64820 10444 64830 10500
rect 65538 10444 65548 10500
rect 65604 10444 67564 10500
rect 67620 10444 67630 10500
rect 31892 10332 35588 10388
rect 47842 10332 47852 10388
rect 47908 10332 48636 10388
rect 48692 10332 48702 10388
rect 54674 10332 54684 10388
rect 54740 10332 56028 10388
rect 56084 10332 56094 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 31892 10164 31948 10332
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 35532 10164 35588 10332
rect 61180 10276 61236 10444
rect 71148 10388 71204 10780
rect 115836 10724 115892 10780
rect 73714 10668 73724 10724
rect 73780 10668 74172 10724
rect 74228 10668 74238 10724
rect 74946 10668 74956 10724
rect 75012 10668 76188 10724
rect 76244 10668 76254 10724
rect 82674 10668 82684 10724
rect 82740 10668 87612 10724
rect 87668 10668 87678 10724
rect 97412 10668 103516 10724
rect 103572 10668 104188 10724
rect 104244 10668 105308 10724
rect 105364 10668 105374 10724
rect 114258 10668 114268 10724
rect 114324 10668 115612 10724
rect 115668 10668 115678 10724
rect 115836 10668 120204 10724
rect 120260 10668 120270 10724
rect 97412 10612 97468 10668
rect 73378 10556 73388 10612
rect 73444 10556 74844 10612
rect 74900 10556 74910 10612
rect 91074 10556 91084 10612
rect 91140 10556 97468 10612
rect 100146 10556 100156 10612
rect 100212 10556 107884 10612
rect 107940 10556 108332 10612
rect 108388 10556 109004 10612
rect 109060 10556 109070 10612
rect 109172 10556 130732 10612
rect 130788 10556 130798 10612
rect 109172 10500 109228 10556
rect 73826 10444 73836 10500
rect 73892 10444 76188 10500
rect 76244 10444 78876 10500
rect 78932 10444 79772 10500
rect 79828 10444 81228 10500
rect 81284 10444 82236 10500
rect 82292 10444 82684 10500
rect 82740 10444 82750 10500
rect 88274 10444 88284 10500
rect 88340 10444 91644 10500
rect 91700 10444 91710 10500
rect 95106 10444 95116 10500
rect 95172 10444 97244 10500
rect 97300 10444 97804 10500
rect 97860 10444 97870 10500
rect 99698 10444 99708 10500
rect 99764 10444 102788 10500
rect 102946 10444 102956 10500
rect 103012 10444 109228 10500
rect 112018 10444 112028 10500
rect 112084 10444 117124 10500
rect 117254 10444 117292 10500
rect 117348 10444 117358 10500
rect 118178 10444 118188 10500
rect 118244 10444 156268 10500
rect 156324 10444 156334 10500
rect 102732 10388 102788 10444
rect 117068 10388 117124 10444
rect 36978 10220 36988 10276
rect 37044 10220 38108 10276
rect 38164 10220 61236 10276
rect 61292 10332 71148 10388
rect 71204 10332 71214 10388
rect 72044 10332 85484 10388
rect 85540 10332 85550 10388
rect 85652 10332 99484 10388
rect 99540 10332 99550 10388
rect 102732 10332 104076 10388
rect 104132 10332 106428 10388
rect 106484 10332 106652 10388
rect 106708 10332 106718 10388
rect 106978 10332 106988 10388
rect 107044 10332 108668 10388
rect 108724 10332 108734 10388
rect 109778 10332 109788 10388
rect 109844 10332 116060 10388
rect 116116 10332 116126 10388
rect 117068 10332 119980 10388
rect 120036 10332 120046 10388
rect 120194 10332 120204 10388
rect 120260 10332 172172 10388
rect 172228 10332 172238 10388
rect 61292 10164 61348 10332
rect 72044 10276 72100 10332
rect 85652 10276 85708 10332
rect 67778 10220 67788 10276
rect 67844 10220 68124 10276
rect 68180 10220 72100 10276
rect 78418 10220 78428 10276
rect 78484 10220 85708 10276
rect 95330 10220 95340 10276
rect 95396 10220 96012 10276
rect 96068 10220 96078 10276
rect 97010 10220 97020 10276
rect 97076 10220 99596 10276
rect 99652 10220 99662 10276
rect 102722 10220 102732 10276
rect 102788 10220 103292 10276
rect 103348 10220 103964 10276
rect 104020 10220 108556 10276
rect 108612 10220 109340 10276
rect 109396 10220 109406 10276
rect 109890 10220 109900 10276
rect 109956 10220 113148 10276
rect 113204 10220 118188 10276
rect 118244 10220 118254 10276
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 96626 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96910 10220
rect 127346 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127630 10220
rect 158066 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158350 10220
rect 18610 10108 18620 10164
rect 18676 10108 31948 10164
rect 35532 10108 61348 10164
rect 62626 10108 62636 10164
rect 62692 10108 63196 10164
rect 63252 10108 63262 10164
rect 64754 10108 64764 10164
rect 64820 10108 65548 10164
rect 65604 10108 65614 10164
rect 71810 10108 71820 10164
rect 71876 10108 75292 10164
rect 75348 10108 75358 10164
rect 87602 10108 87612 10164
rect 87668 10108 88284 10164
rect 88340 10108 88956 10164
rect 89012 10108 89022 10164
rect 98690 10108 98700 10164
rect 98756 10108 103068 10164
rect 103124 10108 105364 10164
rect 105522 10108 105532 10164
rect 105588 10108 106092 10164
rect 106148 10108 113428 10164
rect 113586 10108 113596 10164
rect 113652 10108 114268 10164
rect 114324 10108 114334 10164
rect 114482 10108 114492 10164
rect 114548 10108 115948 10164
rect 116004 10108 116014 10164
rect 128482 10108 128492 10164
rect 128548 10108 129052 10164
rect 129108 10108 135660 10164
rect 135716 10108 135726 10164
rect 105308 10052 105364 10108
rect 113372 10052 113428 10108
rect 36306 9996 36316 10052
rect 36372 9996 39900 10052
rect 39956 9996 39966 10052
rect 49074 9996 49084 10052
rect 49140 9996 51212 10052
rect 51268 9996 52332 10052
rect 52388 9996 52398 10052
rect 71250 9996 71260 10052
rect 71316 9996 71932 10052
rect 71988 9996 71998 10052
rect 81666 9996 81676 10052
rect 81732 9996 83580 10052
rect 83636 9996 83646 10052
rect 85250 9996 85260 10052
rect 85316 9996 85820 10052
rect 85876 9996 85886 10052
rect 87490 9996 87500 10052
rect 87556 9996 88172 10052
rect 88228 9996 88238 10052
rect 95554 9996 95564 10052
rect 95620 9996 96348 10052
rect 96404 9996 96414 10052
rect 105308 9996 106764 10052
rect 106820 9996 112140 10052
rect 112196 9996 112206 10052
rect 113372 9996 114996 10052
rect 116386 9996 116396 10052
rect 116452 9996 119308 10052
rect 119364 9996 119374 10052
rect 53666 9884 53676 9940
rect 53732 9884 53900 9940
rect 53956 9884 55020 9940
rect 55076 9884 55086 9940
rect 62290 9884 62300 9940
rect 62356 9884 63420 9940
rect 63476 9884 65772 9940
rect 65828 9884 66556 9940
rect 66612 9884 66622 9940
rect 84466 9884 84476 9940
rect 84532 9884 84588 9940
rect 84644 9884 84654 9940
rect 111794 9884 111804 9940
rect 111860 9884 114156 9940
rect 114212 9884 114222 9940
rect 66556 9828 66612 9884
rect 114940 9828 114996 9996
rect 115154 9884 115164 9940
rect 115220 9884 125244 9940
rect 125300 9884 125310 9940
rect 66556 9772 68348 9828
rect 68404 9772 68796 9828
rect 68852 9772 68862 9828
rect 77186 9772 77196 9828
rect 77252 9772 77756 9828
rect 77812 9772 81004 9828
rect 81060 9772 81452 9828
rect 81508 9772 81788 9828
rect 81844 9772 82236 9828
rect 82292 9772 82302 9828
rect 99138 9772 99148 9828
rect 99204 9772 100268 9828
rect 100324 9772 100334 9828
rect 113894 9772 113932 9828
rect 113988 9772 113998 9828
rect 114940 9772 119756 9828
rect 119812 9772 119822 9828
rect 36530 9660 36540 9716
rect 36596 9660 51548 9716
rect 51604 9660 51614 9716
rect 74722 9660 74732 9716
rect 74788 9660 75180 9716
rect 75236 9660 75246 9716
rect 78754 9660 78764 9716
rect 78820 9660 79212 9716
rect 79268 9660 84924 9716
rect 84980 9660 84990 9716
rect 87602 9660 87612 9716
rect 87668 9660 89068 9716
rect 89124 9660 89134 9716
rect 93986 9660 93996 9716
rect 94052 9660 96572 9716
rect 96628 9660 96638 9716
rect 98354 9660 98364 9716
rect 98420 9660 98812 9716
rect 98868 9660 98878 9716
rect 112130 9660 112140 9716
rect 112196 9660 114492 9716
rect 114548 9660 114558 9716
rect 116610 9660 116620 9716
rect 116676 9660 117292 9716
rect 117348 9660 118412 9716
rect 118468 9660 119196 9716
rect 119252 9660 119262 9716
rect 30706 9548 30716 9604
rect 30772 9548 32844 9604
rect 32900 9548 33964 9604
rect 34020 9548 37660 9604
rect 37716 9548 37726 9604
rect 43652 9548 55468 9604
rect 55682 9548 55692 9604
rect 55748 9548 56364 9604
rect 56420 9548 56430 9604
rect 62514 9548 62524 9604
rect 62580 9548 62972 9604
rect 63028 9548 65212 9604
rect 65268 9548 65436 9604
rect 65492 9548 65502 9604
rect 73892 9548 80108 9604
rect 80164 9548 82348 9604
rect 82404 9548 82908 9604
rect 82964 9548 82974 9604
rect 83122 9548 83132 9604
rect 83188 9548 85148 9604
rect 85204 9548 85214 9604
rect 94994 9548 95004 9604
rect 95060 9548 97468 9604
rect 97524 9548 97534 9604
rect 97682 9548 97692 9604
rect 97748 9548 99372 9604
rect 99428 9548 99820 9604
rect 99876 9548 100380 9604
rect 100436 9548 100940 9604
rect 100996 9548 101276 9604
rect 101332 9548 101342 9604
rect 104178 9548 104188 9604
rect 104244 9548 105980 9604
rect 106036 9548 106046 9604
rect 110002 9548 110012 9604
rect 110068 9548 112812 9604
rect 112868 9548 118636 9604
rect 118692 9548 118702 9604
rect 39890 9436 39900 9492
rect 39956 9436 43484 9492
rect 43540 9436 43550 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 43652 9380 43708 9548
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 55412 9380 55468 9548
rect 73892 9492 73948 9548
rect 98364 9492 98420 9548
rect 68562 9436 68572 9492
rect 68628 9436 68796 9492
rect 68852 9436 73948 9492
rect 75282 9436 75292 9492
rect 75348 9436 76860 9492
rect 76916 9436 79660 9492
rect 79716 9436 81004 9492
rect 81060 9436 81070 9492
rect 82562 9436 82572 9492
rect 82628 9436 83692 9492
rect 83748 9436 86156 9492
rect 86212 9436 87500 9492
rect 87556 9436 87566 9492
rect 98354 9436 98364 9492
rect 98420 9436 98430 9492
rect 81266 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81550 9436
rect 111986 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112270 9436
rect 142706 9380 142716 9436
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142980 9380 142990 9436
rect 173426 9380 173436 9436
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173700 9380 173710 9436
rect 22754 9324 22764 9380
rect 22820 9324 43708 9380
rect 45714 9324 45724 9380
rect 45780 9324 46172 9380
rect 46228 9324 46238 9380
rect 55412 9324 72716 9380
rect 72772 9324 73276 9380
rect 73332 9324 73342 9380
rect 97794 9324 97804 9380
rect 97860 9324 99148 9380
rect 99204 9324 99214 9380
rect 115490 9324 115500 9380
rect 115556 9324 115948 9380
rect 116004 9324 116014 9380
rect 40114 9212 40124 9268
rect 40180 9212 41916 9268
rect 41972 9212 41982 9268
rect 45826 9212 45836 9268
rect 45892 9212 45902 9268
rect 46834 9212 46844 9268
rect 46900 9212 48972 9268
rect 49028 9212 49038 9268
rect 55010 9212 55020 9268
rect 55076 9212 63868 9268
rect 63924 9212 64204 9268
rect 64260 9212 64270 9268
rect 65426 9212 65436 9268
rect 65492 9212 66220 9268
rect 66276 9212 66892 9268
rect 66948 9212 67788 9268
rect 67844 9212 68684 9268
rect 68740 9212 68750 9268
rect 73714 9212 73724 9268
rect 73780 9212 75404 9268
rect 75460 9212 76300 9268
rect 76356 9212 77532 9268
rect 77588 9212 78540 9268
rect 78596 9212 78606 9268
rect 79650 9212 79660 9268
rect 79716 9212 80444 9268
rect 80500 9212 80780 9268
rect 80836 9212 80846 9268
rect 81554 9212 81564 9268
rect 81620 9212 82572 9268
rect 82628 9212 82638 9268
rect 90178 9212 90188 9268
rect 90244 9212 94444 9268
rect 94500 9212 94510 9268
rect 96226 9212 96236 9268
rect 96292 9212 97580 9268
rect 97636 9212 97646 9268
rect 33506 9100 33516 9156
rect 33572 9100 34636 9156
rect 34692 9100 34702 9156
rect 32162 8988 32172 9044
rect 32228 8988 33740 9044
rect 33796 8988 33806 9044
rect 34066 8988 34076 9044
rect 34132 8988 35420 9044
rect 35476 8988 35486 9044
rect 37650 8988 37660 9044
rect 37716 8988 37996 9044
rect 38052 8988 41468 9044
rect 41524 8988 41534 9044
rect 43474 8988 43484 9044
rect 43540 8988 43932 9044
rect 43988 8988 44380 9044
rect 44436 8988 44446 9044
rect 35074 8876 35084 8932
rect 35140 8876 35868 8932
rect 35924 8876 35934 8932
rect 38658 8876 38668 8932
rect 38724 8876 39228 8932
rect 39284 8876 39294 8932
rect 45836 8820 45892 9212
rect 97804 9156 97860 9324
rect 100930 9212 100940 9268
rect 100996 9212 114380 9268
rect 114436 9212 114940 9268
rect 114996 9212 115836 9268
rect 115892 9212 115902 9268
rect 120306 9212 120316 9268
rect 120372 9212 120876 9268
rect 120932 9212 120942 9268
rect 121202 9212 121212 9268
rect 121268 9212 121884 9268
rect 121940 9212 121950 9268
rect 46498 9100 46508 9156
rect 46564 9100 47180 9156
rect 47236 9100 47246 9156
rect 48290 9100 48300 9156
rect 48356 9100 48636 9156
rect 48692 9100 49532 9156
rect 49588 9100 49598 9156
rect 55234 9100 55244 9156
rect 55300 9100 55468 9156
rect 55524 9100 56196 9156
rect 58482 9100 58492 9156
rect 58548 9100 58828 9156
rect 58884 9100 59052 9156
rect 59108 9100 59118 9156
rect 59602 9100 59612 9156
rect 59668 9100 61628 9156
rect 61684 9100 61694 9156
rect 65314 9100 65324 9156
rect 65380 9100 78428 9156
rect 78484 9100 78494 9156
rect 85698 9100 85708 9156
rect 85764 9100 88172 9156
rect 88228 9100 88238 9156
rect 94210 9100 94220 9156
rect 94276 9100 97132 9156
rect 97188 9100 97198 9156
rect 97346 9100 97356 9156
rect 97412 9100 98252 9156
rect 98308 9100 98318 9156
rect 99474 9100 99484 9156
rect 99540 9100 99932 9156
rect 99988 9100 100604 9156
rect 100660 9100 100670 9156
rect 108658 9100 108668 9156
rect 108724 9100 113036 9156
rect 113092 9100 113102 9156
rect 116386 9100 116396 9156
rect 116452 9100 117180 9156
rect 117236 9100 117246 9156
rect 117506 9100 117516 9156
rect 117572 9100 119308 9156
rect 119364 9100 119374 9156
rect 56140 9044 56196 9100
rect 49970 8988 49980 9044
rect 50036 8988 50316 9044
rect 50372 8988 53900 9044
rect 53956 8988 53966 9044
rect 54786 8988 54796 9044
rect 54852 8988 55692 9044
rect 55748 8988 55758 9044
rect 56130 8988 56140 9044
rect 56196 8988 56700 9044
rect 56756 8988 58604 9044
rect 58660 8988 58670 9044
rect 59612 8932 59668 9100
rect 60610 8988 60620 9044
rect 60676 8988 61180 9044
rect 61236 8988 62300 9044
rect 62356 8988 62366 9044
rect 62514 8988 62524 9044
rect 62580 8988 62590 9044
rect 63410 8988 63420 9044
rect 63476 8988 64428 9044
rect 64484 8988 64494 9044
rect 69010 8988 69020 9044
rect 69076 8988 72492 9044
rect 72548 8988 72558 9044
rect 74050 8988 74060 9044
rect 74116 8988 74620 9044
rect 74676 8988 74686 9044
rect 75394 8988 75404 9044
rect 75460 8988 83020 9044
rect 83076 8988 86492 9044
rect 86548 8988 101388 9044
rect 101444 8988 102844 9044
rect 102900 8988 104300 9044
rect 104356 8988 107884 9044
rect 107940 8988 109116 9044
rect 109172 8988 109182 9044
rect 110002 8988 110012 9044
rect 110068 8988 112028 9044
rect 112084 8988 115500 9044
rect 115556 8988 115566 9044
rect 120978 8988 120988 9044
rect 121044 8988 121548 9044
rect 121604 8988 148876 9044
rect 148932 8988 148942 9044
rect 58258 8876 58268 8932
rect 58324 8876 59668 8932
rect 31892 8764 43708 8820
rect 45714 8764 45724 8820
rect 45780 8764 52444 8820
rect 52500 8764 52780 8820
rect 52836 8764 53340 8820
rect 53396 8764 53406 8820
rect 31892 8708 31948 8764
rect 15810 8652 15820 8708
rect 15876 8652 31948 8708
rect 43652 8708 43708 8764
rect 62524 8708 62580 8988
rect 62850 8876 62860 8932
rect 62916 8876 64204 8932
rect 64260 8876 64270 8932
rect 67666 8876 67676 8932
rect 67732 8876 68572 8932
rect 68628 8876 68638 8932
rect 69682 8876 69692 8932
rect 69748 8876 72268 8932
rect 72324 8876 72334 8932
rect 77420 8876 78204 8932
rect 78260 8876 78764 8932
rect 78820 8876 78830 8932
rect 80098 8876 80108 8932
rect 80164 8876 80780 8932
rect 80836 8876 80846 8932
rect 81004 8876 83580 8932
rect 83636 8876 83646 8932
rect 88498 8876 88508 8932
rect 88564 8876 93212 8932
rect 93268 8876 104524 8932
rect 104580 8876 105196 8932
rect 105252 8876 105532 8932
rect 105588 8876 105598 8932
rect 109890 8876 109900 8932
rect 109956 8876 115836 8932
rect 115892 8876 115902 8932
rect 117954 8876 117964 8932
rect 118020 8876 119196 8932
rect 119252 8876 119262 8932
rect 123442 8876 123452 8932
rect 123508 8876 139132 8932
rect 139188 8876 139198 8932
rect 69692 8820 69748 8876
rect 77420 8820 77476 8876
rect 81004 8820 81060 8876
rect 64642 8764 64652 8820
rect 64708 8764 69748 8820
rect 77410 8764 77420 8820
rect 77476 8764 77486 8820
rect 80546 8764 80556 8820
rect 80612 8764 81060 8820
rect 82114 8764 82124 8820
rect 82180 8764 84252 8820
rect 84308 8764 84318 8820
rect 96562 8764 96572 8820
rect 96628 8764 99708 8820
rect 99764 8764 99774 8820
rect 105634 8764 105644 8820
rect 105700 8764 108108 8820
rect 108164 8764 110236 8820
rect 110292 8764 110302 8820
rect 113708 8764 124124 8820
rect 124180 8764 124190 8820
rect 124348 8764 140476 8820
rect 140532 8764 140542 8820
rect 113708 8708 113764 8764
rect 124348 8708 124404 8764
rect 43652 8652 62580 8708
rect 68226 8652 68236 8708
rect 68292 8652 68796 8708
rect 68852 8652 68862 8708
rect 78278 8652 78316 8708
rect 78372 8652 78382 8708
rect 81890 8652 81900 8708
rect 81956 8652 82572 8708
rect 82628 8652 82638 8708
rect 100482 8652 100492 8708
rect 100548 8652 101612 8708
rect 101668 8652 101678 8708
rect 102162 8652 102172 8708
rect 102228 8652 109228 8708
rect 109666 8652 109676 8708
rect 109732 8652 113708 8708
rect 113764 8652 113774 8708
rect 114034 8652 114044 8708
rect 114100 8652 114716 8708
rect 114772 8652 114782 8708
rect 116722 8652 116732 8708
rect 116788 8652 117404 8708
rect 117460 8652 117470 8708
rect 119186 8652 119196 8708
rect 119252 8652 119868 8708
rect 119924 8652 119934 8708
rect 124226 8652 124236 8708
rect 124292 8652 124404 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 96626 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96910 8652
rect 109172 8596 109228 8652
rect 127346 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127630 8652
rect 158066 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158350 8652
rect 38994 8540 39004 8596
rect 39060 8540 40236 8596
rect 40292 8540 40302 8596
rect 41346 8540 41356 8596
rect 41412 8540 43036 8596
rect 43092 8540 44828 8596
rect 44884 8540 45500 8596
rect 45556 8540 45566 8596
rect 70018 8540 70028 8596
rect 70084 8540 70812 8596
rect 70868 8540 70878 8596
rect 80098 8540 80108 8596
rect 80164 8540 80668 8596
rect 80724 8540 85036 8596
rect 85092 8540 85102 8596
rect 89618 8540 89628 8596
rect 89684 8540 90300 8596
rect 90356 8540 90366 8596
rect 91858 8540 91868 8596
rect 91924 8540 92428 8596
rect 92484 8540 92494 8596
rect 105186 8540 105196 8596
rect 105252 8540 105980 8596
rect 106036 8540 106046 8596
rect 109172 8540 109564 8596
rect 109620 8540 110796 8596
rect 110852 8540 110862 8596
rect 117282 8540 117292 8596
rect 117348 8540 120148 8596
rect 136770 8540 136780 8596
rect 136836 8540 137788 8596
rect 137844 8540 137854 8596
rect 120092 8484 120148 8540
rect 5954 8428 5964 8484
rect 6020 8428 59276 8484
rect 59332 8428 59342 8484
rect 62178 8428 62188 8484
rect 62244 8428 63756 8484
rect 63812 8428 73836 8484
rect 73892 8428 75404 8484
rect 75460 8428 75470 8484
rect 80434 8428 80444 8484
rect 80500 8428 81620 8484
rect 81778 8428 81788 8484
rect 81844 8428 92988 8484
rect 93044 8428 93772 8484
rect 93828 8428 94108 8484
rect 94164 8428 94174 8484
rect 94770 8428 94780 8484
rect 94836 8428 95228 8484
rect 95284 8428 95294 8484
rect 95666 8428 95676 8484
rect 95732 8428 101276 8484
rect 101332 8428 102396 8484
rect 102452 8428 102462 8484
rect 106082 8428 106092 8484
rect 106148 8428 110012 8484
rect 110068 8428 110078 8484
rect 114482 8428 114492 8484
rect 114548 8428 117964 8484
rect 118020 8428 118030 8484
rect 120092 8428 121044 8484
rect 123890 8428 123900 8484
rect 123956 8428 151340 8484
rect 151396 8428 151406 8484
rect 81564 8372 81620 8428
rect 120988 8372 121044 8428
rect 27794 8316 27804 8372
rect 27860 8316 75292 8372
rect 75348 8316 75358 8372
rect 75506 8316 75516 8372
rect 75572 8316 75852 8372
rect 75908 8316 75918 8372
rect 78530 8316 78540 8372
rect 78596 8316 80668 8372
rect 80724 8316 80734 8372
rect 81564 8316 81676 8372
rect 81732 8316 81742 8372
rect 82114 8316 82124 8372
rect 82180 8316 83692 8372
rect 83748 8316 84812 8372
rect 84868 8316 85820 8372
rect 85876 8316 86268 8372
rect 86324 8316 86334 8372
rect 86930 8316 86940 8372
rect 86996 8316 91644 8372
rect 91700 8316 92428 8372
rect 92484 8316 92494 8372
rect 94210 8316 94220 8372
rect 94276 8316 95340 8372
rect 95396 8316 95788 8372
rect 95844 8316 96684 8372
rect 96740 8316 97244 8372
rect 97300 8316 100156 8372
rect 100212 8316 100222 8372
rect 100380 8316 102396 8372
rect 102452 8316 102462 8372
rect 108434 8316 108444 8372
rect 108500 8316 108780 8372
rect 108836 8316 113260 8372
rect 113316 8316 113326 8372
rect 115714 8316 115724 8372
rect 115780 8316 117180 8372
rect 117236 8316 117246 8372
rect 118738 8316 118748 8372
rect 118804 8316 119980 8372
rect 120036 8316 120046 8372
rect 120978 8316 120988 8372
rect 121044 8316 121054 8372
rect 86268 8260 86324 8316
rect 92428 8260 92484 8316
rect 100380 8260 100436 8316
rect 35074 8204 35084 8260
rect 35140 8204 43708 8260
rect 44034 8204 44044 8260
rect 44100 8204 45724 8260
rect 45780 8204 45790 8260
rect 52546 8204 52556 8260
rect 52612 8204 54012 8260
rect 54068 8204 54078 8260
rect 59266 8204 59276 8260
rect 59332 8204 61404 8260
rect 61460 8204 61470 8260
rect 61628 8204 73948 8260
rect 74498 8204 74508 8260
rect 74564 8204 78988 8260
rect 79044 8204 79054 8260
rect 80882 8204 80892 8260
rect 80948 8204 82012 8260
rect 82068 8204 82078 8260
rect 84700 8204 85484 8260
rect 85540 8204 85550 8260
rect 86268 8204 86828 8260
rect 86884 8204 87276 8260
rect 87332 8204 87342 8260
rect 89506 8204 89516 8260
rect 89572 8204 90188 8260
rect 90244 8204 90254 8260
rect 92428 8204 95452 8260
rect 95508 8204 95518 8260
rect 96338 8204 96348 8260
rect 96404 8204 99148 8260
rect 99204 8204 99214 8260
rect 99372 8204 99708 8260
rect 99764 8204 100436 8260
rect 100594 8204 100604 8260
rect 100660 8204 101388 8260
rect 101444 8204 104412 8260
rect 104468 8204 104860 8260
rect 104916 8204 104926 8260
rect 105522 8204 105532 8260
rect 105588 8204 109340 8260
rect 109396 8204 109406 8260
rect 114706 8204 114716 8260
rect 114772 8204 115164 8260
rect 115220 8204 115230 8260
rect 116050 8204 116060 8260
rect 116116 8204 116956 8260
rect 117012 8204 117022 8260
rect 119074 8204 119084 8260
rect 119140 8204 119644 8260
rect 119700 8204 120652 8260
rect 120708 8204 120718 8260
rect 136630 8204 136668 8260
rect 136724 8204 136734 8260
rect 43652 8148 43708 8204
rect 61628 8148 61684 8204
rect 36418 8092 36428 8148
rect 36484 8092 37324 8148
rect 37380 8092 37390 8148
rect 38882 8092 38892 8148
rect 38948 8092 40348 8148
rect 40404 8092 40414 8148
rect 43652 8092 61684 8148
rect 63858 8092 63868 8148
rect 63924 8092 66444 8148
rect 66500 8092 66510 8148
rect 69458 8092 69468 8148
rect 69524 8092 71260 8148
rect 71316 8092 71326 8148
rect 36866 7980 36876 8036
rect 36932 7980 37772 8036
rect 37828 7980 37838 8036
rect 38892 7924 38948 8092
rect 73892 8036 73948 8204
rect 84700 8148 84756 8204
rect 99372 8148 99428 8204
rect 76514 8092 76524 8148
rect 76580 8092 78540 8148
rect 78596 8092 78606 8148
rect 79874 8092 79884 8148
rect 79940 8092 80556 8148
rect 80612 8092 81340 8148
rect 81396 8092 81406 8148
rect 84690 8092 84700 8148
rect 84756 8092 84766 8148
rect 85026 8092 85036 8148
rect 85092 8092 86492 8148
rect 86548 8092 86716 8148
rect 86772 8092 87500 8148
rect 87556 8092 87566 8148
rect 87826 8092 87836 8148
rect 87892 8092 89292 8148
rect 89348 8092 89358 8148
rect 91970 8092 91980 8148
rect 92036 8092 93100 8148
rect 93156 8092 93166 8148
rect 94546 8092 94556 8148
rect 94612 8092 95004 8148
rect 95060 8092 95070 8148
rect 99250 8092 99260 8148
rect 99316 8092 99428 8148
rect 99810 8092 99820 8148
rect 99876 8092 101612 8148
rect 101668 8092 101678 8148
rect 106866 8092 106876 8148
rect 106932 8092 107212 8148
rect 107268 8092 107278 8148
rect 109452 8092 112252 8148
rect 112308 8092 113708 8148
rect 113764 8092 116508 8148
rect 116564 8092 116574 8148
rect 116722 8092 116732 8148
rect 116788 8092 118076 8148
rect 118132 8092 118142 8148
rect 121202 8092 121212 8148
rect 121268 8092 124236 8148
rect 124292 8092 124302 8148
rect 138898 8092 138908 8148
rect 138964 8092 159068 8148
rect 159124 8092 159134 8148
rect 42242 7980 42252 8036
rect 42308 7980 45052 8036
rect 45108 7980 45118 8036
rect 45714 7980 45724 8036
rect 45780 7980 46396 8036
rect 46452 7980 46462 8036
rect 51874 7980 51884 8036
rect 51940 7980 52332 8036
rect 52388 7980 52398 8036
rect 54226 7980 54236 8036
rect 54292 7980 55916 8036
rect 55972 7980 55982 8036
rect 58370 7980 58380 8036
rect 58436 7980 58716 8036
rect 58772 7980 58782 8036
rect 58930 7980 58940 8036
rect 58996 7980 61516 8036
rect 61572 7980 61582 8036
rect 73892 7980 77868 8036
rect 77924 7980 77934 8036
rect 85250 7980 85260 8036
rect 85316 7980 86940 8036
rect 86996 7980 87006 8036
rect 89394 7980 89404 8036
rect 89460 7980 89852 8036
rect 89908 7980 90860 8036
rect 90916 7980 91308 8036
rect 91364 7980 91374 8036
rect 94770 7980 94780 8036
rect 94836 7980 95564 8036
rect 95620 7980 96236 8036
rect 96292 7980 96302 8036
rect 100146 7980 100156 8036
rect 100212 7980 100828 8036
rect 100884 7980 100894 8036
rect 102358 7980 102396 8036
rect 102452 7980 102462 8036
rect 103506 7980 103516 8036
rect 103572 7980 105084 8036
rect 105140 7980 105756 8036
rect 105812 7980 106652 8036
rect 106708 7980 107996 8036
rect 108052 7980 109228 8036
rect 109284 7980 109294 8036
rect 58716 7924 58772 7980
rect 34514 7868 34524 7924
rect 34580 7868 34748 7924
rect 34804 7868 38948 7924
rect 42578 7868 42588 7924
rect 42644 7868 43036 7924
rect 43092 7868 43102 7924
rect 47282 7868 47292 7924
rect 47348 7868 47358 7924
rect 50978 7868 50988 7924
rect 51044 7868 52220 7924
rect 52276 7868 52286 7924
rect 58716 7868 62300 7924
rect 62356 7868 63756 7924
rect 63812 7868 63822 7924
rect 77522 7868 77532 7924
rect 77588 7868 78876 7924
rect 78932 7868 79212 7924
rect 79268 7868 79278 7924
rect 94882 7868 94892 7924
rect 94948 7868 96124 7924
rect 96180 7868 96460 7924
rect 96516 7868 96526 7924
rect 97346 7868 97356 7924
rect 97412 7868 97580 7924
rect 97636 7868 97646 7924
rect 97794 7868 97804 7924
rect 97860 7868 98252 7924
rect 98308 7868 100996 7924
rect 101490 7868 101500 7924
rect 101556 7868 102956 7924
rect 103012 7868 106876 7924
rect 106932 7868 107884 7924
rect 107940 7868 107950 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 43036 7812 43092 7868
rect 47292 7812 47348 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 81266 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81550 7868
rect 26786 7756 26796 7812
rect 26852 7756 27804 7812
rect 27860 7756 27870 7812
rect 43036 7756 43708 7812
rect 43764 7756 43774 7812
rect 43922 7756 43932 7812
rect 43988 7756 44828 7812
rect 44884 7756 47348 7812
rect 55412 7756 75516 7812
rect 75572 7756 75582 7812
rect 75730 7756 75740 7812
rect 75796 7756 76524 7812
rect 76580 7756 76590 7812
rect 77746 7756 77756 7812
rect 77812 7756 78428 7812
rect 78484 7756 78494 7812
rect 95218 7756 95228 7812
rect 95284 7756 97692 7812
rect 97748 7756 97758 7812
rect 99586 7756 99596 7812
rect 99652 7756 100492 7812
rect 100548 7756 100558 7812
rect 55412 7700 55468 7756
rect 100940 7700 100996 7868
rect 109452 7812 109508 8092
rect 111122 7980 111132 8036
rect 111188 7980 112588 8036
rect 112644 7980 114156 8036
rect 114212 7980 114828 8036
rect 114884 7980 114894 8036
rect 115714 7980 115724 8036
rect 115780 7980 118300 8036
rect 118356 7980 118366 8036
rect 118738 7980 118748 8036
rect 118804 7980 119756 8036
rect 119812 7980 119822 8036
rect 120418 7980 120428 8036
rect 120484 7980 120764 8036
rect 120820 7980 121996 8036
rect 122052 7980 122062 8036
rect 130162 7980 130172 8036
rect 130228 7980 130620 8036
rect 130676 7980 130686 8036
rect 131058 7980 131068 8036
rect 131124 7980 171276 8036
rect 171332 7980 171342 8036
rect 130620 7924 130676 7980
rect 112802 7868 112812 7924
rect 112868 7868 116172 7924
rect 116228 7868 116238 7924
rect 118850 7868 118860 7924
rect 118916 7868 121884 7924
rect 121940 7868 121950 7924
rect 130620 7868 142548 7924
rect 111986 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112270 7868
rect 107650 7756 107660 7812
rect 107716 7756 109508 7812
rect 110012 7756 111692 7812
rect 111748 7756 111758 7812
rect 112354 7756 112364 7812
rect 112420 7756 118412 7812
rect 118468 7756 119532 7812
rect 119588 7756 119598 7812
rect 120932 7756 122220 7812
rect 122276 7756 122286 7812
rect 135538 7756 135548 7812
rect 135604 7756 138012 7812
rect 138068 7756 138078 7812
rect 110012 7700 110068 7756
rect 120932 7700 120988 7756
rect 142492 7700 142548 7868
rect 142706 7812 142716 7868
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142980 7812 142990 7868
rect 173426 7812 173436 7868
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173700 7812 173710 7868
rect 29138 7644 29148 7700
rect 29204 7644 55468 7700
rect 57026 7644 57036 7700
rect 57092 7644 57484 7700
rect 57540 7644 59164 7700
rect 59220 7644 59230 7700
rect 61282 7644 61292 7700
rect 61348 7644 62412 7700
rect 62468 7644 62478 7700
rect 75394 7644 75404 7700
rect 75460 7644 79772 7700
rect 79828 7644 79838 7700
rect 80770 7644 80780 7700
rect 80836 7644 81564 7700
rect 81620 7644 93548 7700
rect 93604 7644 93614 7700
rect 94406 7644 94444 7700
rect 94500 7644 95340 7700
rect 95396 7644 96068 7700
rect 97010 7644 97020 7700
rect 97076 7644 97244 7700
rect 97300 7644 98028 7700
rect 98084 7644 99708 7700
rect 99764 7644 99774 7700
rect 100930 7644 100940 7700
rect 100996 7644 101500 7700
rect 101556 7644 105532 7700
rect 105588 7644 105598 7700
rect 107090 7644 107100 7700
rect 107156 7644 107436 7700
rect 107492 7644 107502 7700
rect 108546 7644 108556 7700
rect 108612 7644 110068 7700
rect 110226 7644 110236 7700
rect 110292 7644 114380 7700
rect 114436 7644 114716 7700
rect 114772 7644 114782 7700
rect 118514 7644 118524 7700
rect 118580 7644 120988 7700
rect 121314 7644 121324 7700
rect 121380 7644 123228 7700
rect 123284 7644 123294 7700
rect 129266 7644 129276 7700
rect 129332 7644 129948 7700
rect 130004 7644 130014 7700
rect 130274 7644 130284 7700
rect 130340 7644 130844 7700
rect 130900 7644 132412 7700
rect 132468 7644 132478 7700
rect 133074 7644 133084 7700
rect 133140 7644 133532 7700
rect 133588 7644 134428 7700
rect 134484 7644 134494 7700
rect 142492 7644 143948 7700
rect 144004 7644 144014 7700
rect 96012 7588 96068 7644
rect 32274 7532 32284 7588
rect 32340 7532 35420 7588
rect 35476 7532 35486 7588
rect 42802 7532 42812 7588
rect 42868 7532 44156 7588
rect 44212 7532 44222 7588
rect 60722 7532 60732 7588
rect 60788 7532 60956 7588
rect 61012 7532 67116 7588
rect 67172 7532 67182 7588
rect 75506 7532 75516 7588
rect 75572 7532 79884 7588
rect 79940 7532 79950 7588
rect 81666 7532 81676 7588
rect 81732 7532 85708 7588
rect 87714 7532 87724 7588
rect 87780 7532 90748 7588
rect 90804 7532 90814 7588
rect 93986 7532 93996 7588
rect 94052 7532 95228 7588
rect 95284 7532 95294 7588
rect 95638 7532 95676 7588
rect 95732 7532 95742 7588
rect 96012 7532 98140 7588
rect 98196 7532 98206 7588
rect 104178 7532 104188 7588
rect 104244 7532 105756 7588
rect 105812 7532 106204 7588
rect 106260 7532 107996 7588
rect 108052 7532 108062 7588
rect 115938 7532 115948 7588
rect 116004 7532 118860 7588
rect 118916 7532 118926 7588
rect 119634 7532 119644 7588
rect 119700 7532 121436 7588
rect 121492 7532 121502 7588
rect 128594 7532 128604 7588
rect 128660 7532 164332 7588
rect 164388 7532 164398 7588
rect 85652 7476 85708 7532
rect 33058 7420 33068 7476
rect 33124 7420 33516 7476
rect 33572 7420 36092 7476
rect 36148 7420 36158 7476
rect 46946 7420 46956 7476
rect 47012 7420 48748 7476
rect 48804 7420 48814 7476
rect 55346 7420 55356 7476
rect 55412 7420 55580 7476
rect 55636 7420 55804 7476
rect 55860 7420 55870 7476
rect 66434 7420 66444 7476
rect 66500 7420 66892 7476
rect 66948 7420 69356 7476
rect 69412 7420 69422 7476
rect 71250 7420 71260 7476
rect 71316 7420 71596 7476
rect 71652 7420 74508 7476
rect 74564 7420 74574 7476
rect 75282 7420 75292 7476
rect 75348 7420 77644 7476
rect 77700 7420 77710 7476
rect 80994 7420 81004 7476
rect 81060 7420 81228 7476
rect 81284 7420 82348 7476
rect 82404 7420 82414 7476
rect 83458 7420 83468 7476
rect 83524 7420 84028 7476
rect 84084 7420 84094 7476
rect 85652 7420 93772 7476
rect 93828 7420 93838 7476
rect 98578 7420 98588 7476
rect 98644 7420 100492 7476
rect 100548 7420 101052 7476
rect 101108 7420 102732 7476
rect 102788 7420 103628 7476
rect 103684 7420 106428 7476
rect 106484 7420 106494 7476
rect 106876 7420 110796 7476
rect 110852 7420 110862 7476
rect 114706 7420 114716 7476
rect 114772 7420 115388 7476
rect 115444 7420 115724 7476
rect 115780 7420 115790 7476
rect 117618 7420 117628 7476
rect 117684 7420 118524 7476
rect 118580 7420 118748 7476
rect 118804 7420 119476 7476
rect 18274 7308 18284 7364
rect 18340 7308 19292 7364
rect 19348 7308 21532 7364
rect 21588 7308 22428 7364
rect 22484 7308 25676 7364
rect 25732 7308 25742 7364
rect 31042 7308 31052 7364
rect 31108 7308 31948 7364
rect 35298 7308 35308 7364
rect 35364 7308 39004 7364
rect 39060 7308 41356 7364
rect 41412 7308 41422 7364
rect 46162 7308 46172 7364
rect 46228 7308 46732 7364
rect 46788 7308 48412 7364
rect 48468 7308 49756 7364
rect 49812 7308 49822 7364
rect 61394 7308 61404 7364
rect 61460 7308 69804 7364
rect 69860 7308 69870 7364
rect 71026 7308 71036 7364
rect 71092 7308 71708 7364
rect 71764 7308 71774 7364
rect 76514 7308 76524 7364
rect 76580 7308 77084 7364
rect 77140 7308 77150 7364
rect 77858 7308 77868 7364
rect 77924 7308 83916 7364
rect 83972 7308 87724 7364
rect 87780 7308 88508 7364
rect 88564 7308 88732 7364
rect 88788 7308 88798 7364
rect 96086 7308 96124 7364
rect 96180 7308 97244 7364
rect 97300 7308 98700 7364
rect 98756 7308 98766 7364
rect 99138 7308 99148 7364
rect 99204 7308 100380 7364
rect 100436 7308 100446 7364
rect 31892 7252 31948 7308
rect 88732 7252 88788 7308
rect 99148 7252 99204 7308
rect 106876 7252 106932 7420
rect 119420 7364 119476 7420
rect 120092 7420 122444 7476
rect 122500 7420 122510 7476
rect 130050 7420 130060 7476
rect 130116 7420 130396 7476
rect 130452 7420 131964 7476
rect 132020 7420 132030 7476
rect 21970 7196 21980 7252
rect 22036 7196 24332 7252
rect 24388 7196 24398 7252
rect 31892 7196 32844 7252
rect 32900 7196 34188 7252
rect 34244 7196 47852 7252
rect 47908 7196 48636 7252
rect 48692 7196 48702 7252
rect 68898 7196 68908 7252
rect 68964 7196 69692 7252
rect 69748 7196 69758 7252
rect 75282 7196 75292 7252
rect 75348 7196 75628 7252
rect 75684 7196 75694 7252
rect 77522 7196 77532 7252
rect 77588 7196 78204 7252
rect 78260 7196 78270 7252
rect 81666 7196 81676 7252
rect 81732 7196 84028 7252
rect 84084 7196 84094 7252
rect 88732 7196 89740 7252
rect 89796 7196 90188 7252
rect 90244 7196 90254 7252
rect 93202 7196 93212 7252
rect 93268 7196 97580 7252
rect 97636 7196 97646 7252
rect 98130 7196 98140 7252
rect 98196 7196 99204 7252
rect 104178 7196 104188 7252
rect 104244 7196 106932 7252
rect 106988 7308 111580 7364
rect 111636 7308 112028 7364
rect 112084 7308 113484 7364
rect 113540 7308 113820 7364
rect 113876 7308 113886 7364
rect 114258 7308 114268 7364
rect 114324 7308 118972 7364
rect 119028 7308 119038 7364
rect 119410 7308 119420 7364
rect 119476 7308 119486 7364
rect 106988 7140 107044 7308
rect 120092 7252 120148 7420
rect 120306 7308 120316 7364
rect 120372 7308 121324 7364
rect 121380 7308 121390 7364
rect 121986 7308 121996 7364
rect 122052 7308 132748 7364
rect 137442 7308 137452 7364
rect 137508 7308 138796 7364
rect 138852 7308 138862 7364
rect 140438 7308 140476 7364
rect 140532 7308 140542 7364
rect 132692 7252 132748 7308
rect 109442 7196 109452 7252
rect 109508 7196 112812 7252
rect 112868 7196 112878 7252
rect 113894 7196 113932 7252
rect 113988 7196 113998 7252
rect 114146 7196 114156 7252
rect 114212 7196 114716 7252
rect 114772 7196 114782 7252
rect 115154 7196 115164 7252
rect 115220 7196 115836 7252
rect 115892 7196 115902 7252
rect 118178 7196 118188 7252
rect 118244 7196 120148 7252
rect 122434 7196 122444 7252
rect 122500 7196 127764 7252
rect 132692 7196 137788 7252
rect 127708 7140 127764 7196
rect 137732 7140 137788 7196
rect 22082 7084 22092 7140
rect 22148 7084 24220 7140
rect 24276 7084 31276 7140
rect 31332 7084 31948 7140
rect 45826 7084 45836 7140
rect 45892 7084 57148 7140
rect 57204 7084 57932 7140
rect 57988 7084 59724 7140
rect 59780 7084 59790 7140
rect 68002 7084 68012 7140
rect 68068 7084 69468 7140
rect 69524 7084 69534 7140
rect 82086 7084 82124 7140
rect 82180 7084 82190 7140
rect 97244 7084 98252 7140
rect 98308 7084 98318 7140
rect 106642 7084 106652 7140
rect 106708 7084 107044 7140
rect 108210 7084 108220 7140
rect 108276 7084 109004 7140
rect 109060 7084 117292 7140
rect 117348 7084 117358 7140
rect 118962 7084 118972 7140
rect 119028 7084 121100 7140
rect 121156 7084 121166 7140
rect 127708 7084 134652 7140
rect 134708 7084 134718 7140
rect 137732 7084 138236 7140
rect 138292 7084 138302 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 31892 6916 31948 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 96626 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96910 7084
rect 97244 7028 97300 7084
rect 127346 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127630 7084
rect 158066 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158350 7084
rect 50418 6972 50428 7028
rect 50484 6972 51212 7028
rect 51268 6972 51278 7028
rect 62962 6972 62972 7028
rect 63028 6972 63532 7028
rect 63588 6972 63598 7028
rect 67172 6972 71260 7028
rect 71316 6972 71326 7028
rect 73892 6972 76412 7028
rect 76468 6972 83020 7028
rect 83076 6972 83086 7028
rect 97234 6972 97244 7028
rect 97300 6972 97310 7028
rect 102386 6972 102396 7028
rect 102452 6972 107100 7028
rect 107156 6972 107166 7028
rect 107986 6972 107996 7028
rect 108052 6972 111244 7028
rect 111300 6972 112364 7028
rect 112420 6972 112430 7028
rect 115154 6972 115164 7028
rect 115220 6972 115500 7028
rect 115556 6972 115566 7028
rect 119522 6972 119532 7028
rect 119588 6972 121772 7028
rect 121828 6972 121838 7028
rect 137302 6972 137340 7028
rect 137396 6972 137406 7028
rect 67172 6916 67228 6972
rect 73892 6916 73948 6972
rect 19954 6860 19964 6916
rect 20020 6860 21980 6916
rect 22036 6860 22046 6916
rect 31892 6860 67228 6916
rect 67788 6860 73948 6916
rect 77298 6860 77308 6916
rect 77364 6860 78092 6916
rect 78148 6860 78158 6916
rect 79426 6860 79436 6916
rect 79492 6860 79772 6916
rect 79828 6860 82236 6916
rect 82292 6860 82302 6916
rect 95218 6860 95228 6916
rect 95284 6860 96236 6916
rect 96292 6860 96302 6916
rect 96674 6860 96684 6916
rect 96740 6860 99260 6916
rect 99316 6860 99326 6916
rect 100146 6860 100156 6916
rect 100212 6860 103964 6916
rect 104020 6860 108556 6916
rect 108612 6860 108622 6916
rect 119298 6860 119308 6916
rect 119364 6860 119868 6916
rect 119924 6860 120092 6916
rect 120148 6860 120158 6916
rect 120428 6860 121996 6916
rect 122052 6860 122062 6916
rect 128930 6860 128940 6916
rect 128996 6860 129006 6916
rect 130946 6860 130956 6916
rect 131012 6860 132300 6916
rect 132356 6860 145180 6916
rect 145236 6860 145246 6916
rect 67788 6804 67844 6860
rect 27794 6748 27804 6804
rect 27860 6748 29148 6804
rect 29204 6748 29214 6804
rect 35970 6748 35980 6804
rect 36036 6748 36540 6804
rect 36596 6748 36606 6804
rect 40898 6748 40908 6804
rect 40964 6748 40974 6804
rect 47618 6748 47628 6804
rect 47684 6748 52108 6804
rect 52164 6748 52174 6804
rect 53778 6748 53788 6804
rect 53844 6748 67844 6804
rect 76178 6748 76188 6804
rect 76244 6748 77532 6804
rect 77588 6748 77598 6804
rect 81218 6748 81228 6804
rect 81284 6748 86380 6804
rect 86436 6748 87276 6804
rect 87332 6748 89852 6804
rect 89908 6748 89918 6804
rect 97682 6748 97692 6804
rect 97748 6748 98588 6804
rect 98644 6748 98654 6804
rect 102498 6748 102508 6804
rect 102564 6748 107212 6804
rect 107268 6748 107278 6804
rect 116060 6748 117404 6804
rect 117460 6748 117852 6804
rect 117908 6748 117918 6804
rect 119074 6748 119084 6804
rect 119140 6748 119756 6804
rect 119812 6748 120204 6804
rect 120260 6748 120270 6804
rect 40908 6692 40964 6748
rect 116060 6692 116116 6748
rect 120428 6692 120484 6860
rect 122098 6748 122108 6804
rect 122164 6748 123452 6804
rect 123508 6748 123518 6804
rect 128146 6748 128156 6804
rect 128212 6748 128604 6804
rect 128660 6748 128670 6804
rect 128940 6692 128996 6860
rect 137526 6748 137564 6804
rect 137620 6748 137630 6804
rect 138226 6748 138236 6804
rect 138292 6748 141260 6804
rect 141316 6748 148988 6804
rect 149044 6748 149054 6804
rect 30594 6636 30604 6692
rect 30660 6636 34860 6692
rect 34916 6636 34926 6692
rect 36418 6636 36428 6692
rect 36484 6636 37436 6692
rect 37492 6636 38220 6692
rect 38276 6636 38286 6692
rect 38770 6636 38780 6692
rect 38836 6636 40628 6692
rect 40908 6636 41804 6692
rect 41860 6636 41870 6692
rect 42466 6636 42476 6692
rect 42532 6636 45612 6692
rect 45668 6636 45678 6692
rect 46162 6636 46172 6692
rect 46228 6636 46396 6692
rect 46452 6636 46462 6692
rect 47730 6636 47740 6692
rect 47796 6636 50876 6692
rect 50932 6636 50942 6692
rect 52210 6636 52220 6692
rect 52276 6636 53452 6692
rect 53508 6636 53518 6692
rect 57110 6636 57148 6692
rect 57204 6636 57214 6692
rect 59714 6636 59724 6692
rect 59780 6636 61852 6692
rect 61908 6636 62300 6692
rect 62356 6636 63420 6692
rect 63476 6636 63486 6692
rect 64866 6636 64876 6692
rect 64932 6636 65660 6692
rect 65716 6636 65726 6692
rect 66098 6636 66108 6692
rect 66164 6636 68124 6692
rect 68180 6636 68190 6692
rect 76626 6636 76636 6692
rect 76692 6636 77308 6692
rect 77364 6636 77374 6692
rect 84466 6636 84476 6692
rect 84532 6636 85260 6692
rect 85316 6636 85326 6692
rect 86706 6636 86716 6692
rect 86772 6636 87500 6692
rect 87556 6636 87566 6692
rect 91494 6636 91532 6692
rect 91588 6636 91598 6692
rect 95106 6636 95116 6692
rect 95172 6636 95900 6692
rect 95956 6636 95966 6692
rect 96226 6636 96236 6692
rect 96292 6636 97468 6692
rect 97524 6636 99484 6692
rect 99540 6636 99932 6692
rect 99988 6636 99998 6692
rect 104150 6636 104188 6692
rect 104244 6636 104254 6692
rect 104402 6636 104412 6692
rect 104468 6636 105084 6692
rect 105140 6636 105150 6692
rect 105298 6636 105308 6692
rect 105364 6636 106092 6692
rect 106148 6636 106158 6692
rect 106726 6636 106764 6692
rect 106820 6636 106830 6692
rect 107090 6636 107100 6692
rect 107156 6636 107324 6692
rect 107380 6636 112140 6692
rect 112196 6636 112206 6692
rect 114034 6636 114044 6692
rect 114100 6636 115948 6692
rect 116004 6636 116116 6692
rect 116610 6636 116620 6692
rect 116676 6636 120484 6692
rect 120642 6636 120652 6692
rect 120708 6636 122444 6692
rect 122500 6636 122780 6692
rect 122836 6636 122846 6692
rect 125682 6636 125692 6692
rect 125748 6636 125916 6692
rect 125972 6636 126924 6692
rect 126980 6636 126990 6692
rect 127820 6636 128996 6692
rect 130610 6636 130620 6692
rect 130676 6636 130844 6692
rect 130900 6636 130910 6692
rect 134754 6636 134764 6692
rect 134820 6636 135884 6692
rect 135940 6636 136892 6692
rect 136948 6636 136958 6692
rect 137330 6636 137340 6692
rect 137396 6636 138684 6692
rect 138740 6636 138750 6692
rect 142034 6636 142044 6692
rect 142100 6636 142716 6692
rect 142772 6636 142782 6692
rect 40572 6580 40628 6636
rect 95900 6580 95956 6636
rect 127820 6580 127876 6636
rect 20178 6524 20188 6580
rect 20244 6524 20636 6580
rect 20692 6524 21532 6580
rect 21588 6524 22540 6580
rect 22596 6524 22876 6580
rect 22932 6524 22942 6580
rect 34178 6524 34188 6580
rect 34244 6524 36204 6580
rect 36260 6524 36270 6580
rect 36642 6524 36652 6580
rect 36708 6524 38892 6580
rect 38948 6524 38958 6580
rect 39666 6524 39676 6580
rect 39732 6524 40348 6580
rect 40404 6524 40414 6580
rect 40562 6524 40572 6580
rect 40628 6524 42140 6580
rect 42196 6524 42206 6580
rect 44034 6524 44044 6580
rect 44100 6524 46284 6580
rect 46340 6524 46508 6580
rect 46564 6524 46574 6580
rect 48962 6524 48972 6580
rect 49028 6524 50148 6580
rect 51314 6524 51324 6580
rect 51380 6524 52332 6580
rect 52388 6524 52398 6580
rect 56578 6524 56588 6580
rect 56644 6524 58044 6580
rect 58100 6524 58110 6580
rect 59378 6524 59388 6580
rect 59444 6524 62636 6580
rect 62692 6524 62702 6580
rect 66770 6524 66780 6580
rect 66836 6524 67676 6580
rect 67732 6524 67742 6580
rect 75954 6524 75964 6580
rect 76020 6524 76524 6580
rect 76580 6524 77756 6580
rect 77812 6524 77822 6580
rect 78306 6524 78316 6580
rect 78372 6524 78428 6580
rect 78484 6524 79772 6580
rect 79828 6524 80444 6580
rect 80500 6524 80510 6580
rect 81442 6524 81452 6580
rect 81508 6524 83916 6580
rect 83972 6524 83982 6580
rect 85810 6524 85820 6580
rect 85876 6524 87052 6580
rect 87108 6524 87118 6580
rect 95900 6524 99036 6580
rect 99092 6524 101836 6580
rect 101892 6524 102620 6580
rect 102676 6524 102686 6580
rect 104514 6524 104524 6580
rect 104580 6524 105644 6580
rect 105700 6524 105710 6580
rect 105858 6524 105868 6580
rect 105924 6524 110348 6580
rect 110404 6524 111188 6580
rect 113026 6524 113036 6580
rect 113092 6524 127820 6580
rect 127876 6524 127886 6580
rect 130060 6524 130508 6580
rect 130564 6524 130574 6580
rect 136658 6524 136668 6580
rect 136724 6524 139132 6580
rect 139188 6524 139804 6580
rect 139860 6524 139870 6580
rect 140130 6524 140140 6580
rect 140196 6524 152572 6580
rect 152628 6524 152638 6580
rect 39676 6468 39732 6524
rect 50092 6468 50148 6524
rect 102620 6468 102676 6524
rect 111132 6468 111188 6524
rect 130060 6468 130116 6524
rect 140140 6468 140196 6524
rect 14914 6412 14924 6468
rect 14980 6412 26068 6468
rect 30930 6412 30940 6468
rect 30996 6412 32060 6468
rect 32116 6412 34972 6468
rect 35028 6412 35038 6468
rect 36866 6412 36876 6468
rect 36932 6412 39732 6468
rect 41794 6412 41804 6468
rect 41860 6412 43820 6468
rect 43876 6412 44604 6468
rect 44660 6412 44670 6468
rect 46386 6412 46396 6468
rect 46452 6412 48188 6468
rect 48244 6412 49644 6468
rect 49700 6412 49710 6468
rect 50092 6412 55244 6468
rect 55300 6412 55310 6468
rect 60386 6412 60396 6468
rect 60452 6412 60844 6468
rect 60900 6412 60910 6468
rect 61730 6412 61740 6468
rect 61796 6412 64316 6468
rect 64372 6412 64382 6468
rect 65762 6412 65772 6468
rect 65828 6412 66556 6468
rect 66612 6412 66622 6468
rect 66994 6412 67004 6468
rect 67060 6412 70028 6468
rect 70084 6412 70094 6468
rect 70914 6412 70924 6468
rect 70980 6412 72044 6468
rect 72100 6412 72110 6468
rect 77410 6412 77420 6468
rect 77476 6412 82348 6468
rect 82404 6412 82414 6468
rect 84130 6412 84140 6468
rect 84196 6412 84588 6468
rect 84644 6412 85484 6468
rect 85540 6412 85550 6468
rect 87826 6412 87836 6468
rect 87892 6412 88172 6468
rect 88228 6412 90524 6468
rect 90580 6412 90590 6468
rect 102620 6412 105980 6468
rect 106036 6412 106046 6468
rect 109330 6412 109340 6468
rect 109396 6412 109564 6468
rect 109620 6412 109630 6468
rect 111122 6412 111132 6468
rect 111188 6412 111198 6468
rect 111356 6412 114268 6468
rect 114324 6412 114334 6468
rect 116274 6412 116284 6468
rect 116340 6412 118748 6468
rect 118804 6412 118814 6468
rect 120082 6412 120092 6468
rect 120148 6412 120988 6468
rect 121986 6412 121996 6468
rect 122052 6412 122780 6468
rect 122836 6412 122846 6468
rect 123890 6412 123900 6468
rect 123956 6412 123966 6468
rect 128034 6412 128044 6468
rect 128100 6412 128492 6468
rect 128548 6412 128558 6468
rect 130050 6412 130060 6468
rect 130116 6412 130126 6468
rect 133858 6412 133868 6468
rect 133924 6412 133934 6468
rect 135762 6412 135772 6468
rect 135828 6412 137228 6468
rect 137284 6412 137788 6468
rect 139346 6412 139356 6468
rect 139412 6412 140196 6468
rect 142370 6412 142380 6468
rect 142436 6412 142604 6468
rect 142660 6412 143052 6468
rect 143108 6412 143118 6468
rect 145730 6412 145740 6468
rect 145796 6412 146636 6468
rect 146692 6412 146972 6468
rect 147028 6412 147038 6468
rect 26012 6356 26068 6412
rect 16370 6300 16380 6356
rect 16436 6300 17388 6356
rect 17444 6300 18844 6356
rect 18900 6300 19180 6356
rect 19236 6300 19246 6356
rect 23202 6300 23212 6356
rect 23268 6300 23548 6356
rect 23604 6300 23614 6356
rect 26012 6300 42028 6356
rect 42084 6300 42700 6356
rect 42756 6300 42766 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 23548 6244 23604 6300
rect 14802 6188 14812 6244
rect 14868 6188 17724 6244
rect 17780 6188 18396 6244
rect 18452 6188 18462 6244
rect 23548 6188 31052 6244
rect 31108 6188 31118 6244
rect 40450 6188 40460 6244
rect 40516 6188 41356 6244
rect 41412 6188 42812 6244
rect 42868 6188 42878 6244
rect 44604 6132 44660 6412
rect 64316 6356 64372 6412
rect 111356 6356 111412 6412
rect 120932 6356 120988 6412
rect 123900 6356 123956 6412
rect 133868 6356 133924 6412
rect 137732 6356 137788 6412
rect 46050 6300 46060 6356
rect 46116 6300 48972 6356
rect 49028 6300 49038 6356
rect 58594 6300 58604 6356
rect 58660 6300 61628 6356
rect 61684 6300 61694 6356
rect 62850 6300 62860 6356
rect 62916 6300 63420 6356
rect 63476 6300 64092 6356
rect 64148 6300 64158 6356
rect 64316 6300 67452 6356
rect 67508 6300 67518 6356
rect 70364 6300 77980 6356
rect 78036 6300 78046 6356
rect 79846 6300 79884 6356
rect 79940 6300 79950 6356
rect 82114 6300 82124 6356
rect 82180 6300 82236 6356
rect 82292 6300 82302 6356
rect 82674 6300 82684 6356
rect 82740 6300 82908 6356
rect 82964 6300 82974 6356
rect 83458 6300 83468 6356
rect 83524 6300 88396 6356
rect 88452 6300 88956 6356
rect 89012 6300 91868 6356
rect 91924 6300 93100 6356
rect 93156 6300 93166 6356
rect 94546 6300 94556 6356
rect 94612 6300 95564 6356
rect 95620 6300 95630 6356
rect 101602 6300 101612 6356
rect 101668 6300 102284 6356
rect 102340 6300 102350 6356
rect 103058 6300 103068 6356
rect 103124 6300 103852 6356
rect 103908 6300 103918 6356
rect 104402 6300 104412 6356
rect 104468 6300 108220 6356
rect 108276 6300 108286 6356
rect 110786 6300 110796 6356
rect 110852 6300 111412 6356
rect 114818 6300 114828 6356
rect 114884 6300 116956 6356
rect 117012 6300 117022 6356
rect 119858 6300 119868 6356
rect 119924 6300 120428 6356
rect 120484 6300 120652 6356
rect 120708 6300 120718 6356
rect 120932 6300 123956 6356
rect 124226 6300 124236 6356
rect 124292 6300 124796 6356
rect 124852 6300 132636 6356
rect 132692 6300 134204 6356
rect 134260 6300 134270 6356
rect 137732 6300 139188 6356
rect 140914 6300 140924 6356
rect 140980 6300 142268 6356
rect 142324 6300 142334 6356
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 62860 6244 62916 6300
rect 70364 6244 70420 6300
rect 81266 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81550 6300
rect 111986 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112270 6300
rect 45938 6188 45948 6244
rect 46004 6188 47628 6244
rect 47684 6188 47694 6244
rect 54786 6188 54796 6244
rect 54852 6188 54862 6244
rect 60610 6188 60620 6244
rect 60676 6188 62916 6244
rect 64306 6188 64316 6244
rect 64372 6188 65212 6244
rect 65268 6188 66108 6244
rect 66164 6188 66174 6244
rect 66546 6188 66556 6244
rect 66612 6188 70420 6244
rect 70578 6188 70588 6244
rect 70644 6188 71932 6244
rect 71988 6188 77756 6244
rect 77812 6188 77822 6244
rect 78866 6188 78876 6244
rect 78932 6188 80780 6244
rect 80836 6188 80846 6244
rect 82450 6188 82460 6244
rect 82516 6188 85596 6244
rect 85652 6188 86828 6244
rect 86884 6188 88732 6244
rect 88788 6188 89180 6244
rect 89236 6188 90076 6244
rect 90132 6188 90636 6244
rect 90692 6188 90702 6244
rect 92530 6188 92540 6244
rect 92596 6188 95004 6244
rect 95060 6188 95070 6244
rect 113362 6188 113372 6244
rect 113428 6188 115052 6244
rect 115108 6188 116396 6244
rect 116452 6188 116462 6244
rect 117516 6188 123788 6244
rect 123844 6188 123854 6244
rect 54796 6132 54852 6188
rect 117516 6132 117572 6188
rect 124236 6132 124292 6300
rect 139132 6244 139188 6300
rect 142706 6244 142716 6300
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142980 6244 142990 6300
rect 173426 6244 173436 6300
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173700 6244 173710 6300
rect 132934 6188 132972 6244
rect 133028 6188 133038 6244
rect 133186 6188 133196 6244
rect 133252 6188 136220 6244
rect 136276 6188 136286 6244
rect 137330 6188 137340 6244
rect 137396 6188 137676 6244
rect 137732 6188 137742 6244
rect 139122 6188 139132 6244
rect 139188 6188 140028 6244
rect 140084 6188 140700 6244
rect 140756 6188 141708 6244
rect 141764 6188 141774 6244
rect 141708 6132 141764 6188
rect 11554 6076 11564 6132
rect 11620 6076 24724 6132
rect 24882 6076 24892 6132
rect 24948 6076 25676 6132
rect 25732 6076 26908 6132
rect 26964 6076 29036 6132
rect 29092 6076 30604 6132
rect 30660 6076 30670 6132
rect 31892 6076 36988 6132
rect 37044 6076 37054 6132
rect 38098 6076 38108 6132
rect 38164 6076 39340 6132
rect 39396 6076 39406 6132
rect 44604 6076 48076 6132
rect 48132 6076 54852 6132
rect 60386 6076 60396 6132
rect 60452 6076 61068 6132
rect 61124 6076 61134 6132
rect 65538 6076 65548 6132
rect 65604 6076 67228 6132
rect 67284 6076 67294 6132
rect 67778 6076 67788 6132
rect 67844 6076 68796 6132
rect 68852 6076 68862 6132
rect 72258 6076 72268 6132
rect 72324 6076 75404 6132
rect 75460 6076 75470 6132
rect 78988 6076 80108 6132
rect 80164 6076 81452 6132
rect 81508 6076 82348 6132
rect 82404 6076 82414 6132
rect 82562 6076 82572 6132
rect 82628 6076 83132 6132
rect 83188 6076 83468 6132
rect 83524 6076 83534 6132
rect 93762 6076 93772 6132
rect 93828 6076 105644 6132
rect 105700 6076 105710 6132
rect 106866 6076 106876 6132
rect 106932 6076 113484 6132
rect 113540 6076 113550 6132
rect 114034 6076 114044 6132
rect 114100 6076 117572 6132
rect 122220 6076 122332 6132
rect 122388 6076 123340 6132
rect 123396 6076 124292 6132
rect 131170 6076 131180 6132
rect 131236 6076 135324 6132
rect 135380 6076 135390 6132
rect 136966 6076 137004 6132
rect 137060 6076 137070 6132
rect 138674 6076 138684 6132
rect 138740 6076 140812 6132
rect 140868 6076 140878 6132
rect 141708 6076 144956 6132
rect 145012 6076 145022 6132
rect 24668 6020 24724 6076
rect 31892 6020 31948 6076
rect 36988 6020 37044 6076
rect 13458 5964 13468 6020
rect 13524 5964 14924 6020
rect 14980 5964 14990 6020
rect 18386 5964 18396 6020
rect 18452 5964 20076 6020
rect 20132 5964 20142 6020
rect 24668 5964 31948 6020
rect 34178 5964 34188 6020
rect 34244 5964 36764 6020
rect 36820 5964 36830 6020
rect 36988 5964 39564 6020
rect 39620 5964 40460 6020
rect 40516 5964 40526 6020
rect 44146 5964 44156 6020
rect 44212 5964 46172 6020
rect 46228 5964 47628 6020
rect 47684 5964 47694 6020
rect 48850 5964 48860 6020
rect 48916 5964 49980 6020
rect 50036 5964 50046 6020
rect 55682 5964 55692 6020
rect 55748 5964 56364 6020
rect 56420 5964 56430 6020
rect 56690 5964 56700 6020
rect 56756 5964 57484 6020
rect 57540 5964 57550 6020
rect 57698 5964 57708 6020
rect 57764 5964 58268 6020
rect 58324 5964 58334 6020
rect 60498 5964 60508 6020
rect 60564 5964 61292 6020
rect 61348 5964 61358 6020
rect 63634 5964 63644 6020
rect 63700 5964 65100 6020
rect 65156 5964 65166 6020
rect 66322 5964 66332 6020
rect 66388 5964 67900 6020
rect 67956 5964 67966 6020
rect 69318 5964 69356 6020
rect 69412 5964 69422 6020
rect 72370 5964 72380 6020
rect 72436 5964 74060 6020
rect 74116 5964 74126 6020
rect 78988 5908 79044 6076
rect 105644 6020 105700 6076
rect 79986 5964 79996 6020
rect 80052 5964 81340 6020
rect 81396 5964 81406 6020
rect 82674 5964 82684 6020
rect 82740 5964 85484 6020
rect 85540 5964 85550 6020
rect 85652 5964 86044 6020
rect 86100 5964 89068 6020
rect 89124 5964 90972 6020
rect 91028 5964 91644 6020
rect 91700 5964 91710 6020
rect 96226 5964 96236 6020
rect 96292 5964 97356 6020
rect 97412 5964 97422 6020
rect 101154 5964 101164 6020
rect 101220 5964 101836 6020
rect 101892 5964 101902 6020
rect 105644 5964 107100 6020
rect 107156 5964 107166 6020
rect 107426 5964 107436 6020
rect 107492 5964 112588 6020
rect 112644 5964 112654 6020
rect 114930 5964 114940 6020
rect 114996 5964 116396 6020
rect 116452 5964 116462 6020
rect 117618 5964 117628 6020
rect 117684 5964 121996 6020
rect 122052 5964 122062 6020
rect 85652 5908 85708 5964
rect 8194 5852 8204 5908
rect 8260 5852 8652 5908
rect 8708 5852 8718 5908
rect 14354 5852 14364 5908
rect 14420 5852 16604 5908
rect 16660 5852 17388 5908
rect 17444 5852 17454 5908
rect 31490 5852 31500 5908
rect 31556 5852 32620 5908
rect 32676 5852 33964 5908
rect 34020 5852 34030 5908
rect 34738 5852 34748 5908
rect 34804 5852 35532 5908
rect 35588 5852 39452 5908
rect 39508 5852 39518 5908
rect 46274 5852 46284 5908
rect 46340 5852 47404 5908
rect 47460 5852 47470 5908
rect 59602 5852 59612 5908
rect 59668 5852 67564 5908
rect 67620 5852 67630 5908
rect 70690 5852 70700 5908
rect 70756 5852 73164 5908
rect 73220 5852 73388 5908
rect 73444 5852 73454 5908
rect 73938 5852 73948 5908
rect 74004 5852 75516 5908
rect 75572 5852 75582 5908
rect 77970 5852 77980 5908
rect 78036 5852 78988 5908
rect 79044 5852 79054 5908
rect 80322 5852 80332 5908
rect 80388 5852 80398 5908
rect 80658 5852 80668 5908
rect 80724 5852 82124 5908
rect 82180 5852 82190 5908
rect 83234 5852 83244 5908
rect 83300 5852 85036 5908
rect 85092 5852 85102 5908
rect 85484 5852 85708 5908
rect 90738 5852 90748 5908
rect 90804 5852 91980 5908
rect 92036 5852 92046 5908
rect 98914 5852 98924 5908
rect 98980 5852 104972 5908
rect 105028 5852 105038 5908
rect 107986 5852 107996 5908
rect 108052 5852 110348 5908
rect 110404 5852 110796 5908
rect 110852 5852 110862 5908
rect 112690 5852 112700 5908
rect 112756 5852 113148 5908
rect 113204 5852 118076 5908
rect 118132 5852 118142 5908
rect 118626 5852 118636 5908
rect 118692 5852 119868 5908
rect 119924 5852 119934 5908
rect 34748 5796 34804 5852
rect 80332 5796 80388 5852
rect 85484 5796 85540 5852
rect 122220 5796 122276 6076
rect 132972 6020 133028 6076
rect 123666 5964 123676 6020
rect 123732 5964 123788 6020
rect 123844 5964 125356 6020
rect 125412 5964 125422 6020
rect 125794 5964 125804 6020
rect 125860 5964 126476 6020
rect 126532 5964 126542 6020
rect 127922 5964 127932 6020
rect 127988 5964 128604 6020
rect 128660 5964 128670 6020
rect 129602 5964 129612 6020
rect 129668 5964 131740 6020
rect 131796 5964 131806 6020
rect 132962 5964 132972 6020
rect 133028 5964 133038 6020
rect 134530 5964 134540 6020
rect 134596 5964 135772 6020
rect 135828 5964 142380 6020
rect 142436 5964 142446 6020
rect 144498 5964 144508 6020
rect 144564 5964 145292 6020
rect 145348 5964 145740 6020
rect 145796 5964 145806 6020
rect 122658 5852 122668 5908
rect 122724 5852 127708 5908
rect 127764 5852 127774 5908
rect 128258 5852 128268 5908
rect 128324 5852 129276 5908
rect 129332 5852 129342 5908
rect 132692 5852 134652 5908
rect 134708 5852 134718 5908
rect 134866 5852 134876 5908
rect 134932 5852 135996 5908
rect 136052 5852 138124 5908
rect 138180 5852 149548 5908
rect 149604 5852 149614 5908
rect 132692 5796 132748 5852
rect 19842 5740 19852 5796
rect 19908 5740 20524 5796
rect 20580 5740 21196 5796
rect 21252 5740 21262 5796
rect 31602 5740 31612 5796
rect 31668 5740 34804 5796
rect 35074 5740 35084 5796
rect 35140 5740 35756 5796
rect 35812 5740 35822 5796
rect 36866 5740 36876 5796
rect 36932 5740 41748 5796
rect 41906 5740 41916 5796
rect 41972 5740 45276 5796
rect 45332 5740 45500 5796
rect 45556 5740 47964 5796
rect 48020 5740 48030 5796
rect 64418 5740 64428 5796
rect 64484 5740 65436 5796
rect 65492 5740 66780 5796
rect 66836 5740 66846 5796
rect 74694 5740 74732 5796
rect 74788 5740 74798 5796
rect 80332 5740 80892 5796
rect 80948 5740 80958 5796
rect 83010 5740 83020 5796
rect 83076 5740 85540 5796
rect 85652 5740 86492 5796
rect 86548 5740 86558 5796
rect 90962 5740 90972 5796
rect 91028 5740 91532 5796
rect 91588 5740 91598 5796
rect 91746 5740 91756 5796
rect 91812 5740 105420 5796
rect 105476 5740 106540 5796
rect 106596 5740 107436 5796
rect 107492 5740 107502 5796
rect 109442 5740 109452 5796
rect 109508 5740 111020 5796
rect 111076 5740 111086 5796
rect 113586 5740 113596 5796
rect 113652 5740 116228 5796
rect 116386 5740 116396 5796
rect 116452 5740 121100 5796
rect 121156 5740 121166 5796
rect 121426 5740 121436 5796
rect 121492 5740 121996 5796
rect 122052 5740 122276 5796
rect 125010 5740 125020 5796
rect 125076 5740 125580 5796
rect 125636 5740 125646 5796
rect 126802 5740 126812 5796
rect 126868 5740 132748 5796
rect 136630 5740 136668 5796
rect 136724 5740 136734 5796
rect 41692 5684 41748 5740
rect 85652 5684 85708 5740
rect 32050 5628 32060 5684
rect 32116 5628 37492 5684
rect 41692 5628 42812 5684
rect 42868 5628 42878 5684
rect 46610 5628 46620 5684
rect 46676 5628 47852 5684
rect 47908 5628 52444 5684
rect 52500 5628 52510 5684
rect 58594 5628 58604 5684
rect 58660 5628 66668 5684
rect 66724 5628 66734 5684
rect 67442 5628 67452 5684
rect 67508 5628 68796 5684
rect 68852 5628 71372 5684
rect 71428 5628 71438 5684
rect 79874 5628 79884 5684
rect 79940 5628 85708 5684
rect 96002 5628 96012 5684
rect 96068 5628 100716 5684
rect 100772 5628 100782 5684
rect 102386 5628 102396 5684
rect 102452 5628 105644 5684
rect 105700 5628 105710 5684
rect 10658 5516 10668 5572
rect 10724 5516 11228 5572
rect 11284 5516 33068 5572
rect 33124 5516 33134 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 37436 5460 37492 5628
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 71372 5460 71428 5628
rect 84130 5516 84140 5572
rect 84196 5516 85148 5572
rect 85204 5516 91868 5572
rect 91924 5516 91934 5572
rect 104066 5516 104076 5572
rect 104132 5516 105196 5572
rect 105252 5516 107660 5572
rect 107716 5516 107726 5572
rect 111122 5516 111132 5572
rect 111188 5516 113820 5572
rect 113876 5516 113886 5572
rect 96626 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96910 5516
rect 116172 5460 116228 5740
rect 126812 5684 126868 5740
rect 137732 5684 137788 5796
rect 137844 5740 140924 5796
rect 140980 5740 140990 5796
rect 143378 5740 143388 5796
rect 143444 5740 143724 5796
rect 143780 5740 143790 5796
rect 145170 5740 145180 5796
rect 145236 5740 147308 5796
rect 147364 5740 147374 5796
rect 117730 5628 117740 5684
rect 117796 5628 118748 5684
rect 118804 5628 119532 5684
rect 119588 5628 119598 5684
rect 123778 5628 123788 5684
rect 123844 5628 126868 5684
rect 127148 5628 132076 5684
rect 132132 5628 132142 5684
rect 132692 5628 133196 5684
rect 133252 5628 133262 5684
rect 133970 5628 133980 5684
rect 134036 5628 134540 5684
rect 134596 5628 134606 5684
rect 135650 5628 135660 5684
rect 135716 5628 137788 5684
rect 139794 5628 139804 5684
rect 139860 5628 140588 5684
rect 140644 5628 140654 5684
rect 142706 5628 142716 5684
rect 142772 5628 143948 5684
rect 144004 5628 146076 5684
rect 146132 5628 159516 5684
rect 159572 5628 159582 5684
rect 118626 5516 118636 5572
rect 118692 5516 119084 5572
rect 119140 5516 121660 5572
rect 121716 5516 121726 5572
rect 122882 5516 122892 5572
rect 122948 5516 125804 5572
rect 125860 5516 125870 5572
rect 127148 5460 127204 5628
rect 132692 5572 132748 5628
rect 127698 5516 127708 5572
rect 127764 5516 132748 5572
rect 134754 5516 134764 5572
rect 134820 5516 142100 5572
rect 143714 5516 143724 5572
rect 143780 5516 144060 5572
rect 144116 5516 144126 5572
rect 127346 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127630 5516
rect 37426 5404 37436 5460
rect 37492 5404 49084 5460
rect 49140 5404 49150 5460
rect 65090 5404 65100 5460
rect 65156 5404 65548 5460
rect 65604 5404 65614 5460
rect 71372 5404 75068 5460
rect 75124 5404 75134 5460
rect 83570 5404 83580 5460
rect 83636 5404 84252 5460
rect 84308 5404 84700 5460
rect 84756 5404 86604 5460
rect 86660 5404 86670 5460
rect 91634 5404 91644 5460
rect 91700 5404 93660 5460
rect 93716 5404 93726 5460
rect 97412 5404 100268 5460
rect 100324 5404 106652 5460
rect 106708 5404 106718 5460
rect 111346 5404 111356 5460
rect 111412 5404 113708 5460
rect 113764 5404 113932 5460
rect 113988 5404 113998 5460
rect 116172 5404 122108 5460
rect 122164 5404 122174 5460
rect 125570 5404 125580 5460
rect 125636 5404 125916 5460
rect 125972 5404 127204 5460
rect 130050 5404 130060 5460
rect 130116 5404 132748 5460
rect 133830 5404 133868 5460
rect 133924 5404 133934 5460
rect 134530 5404 134540 5460
rect 134596 5404 135548 5460
rect 135604 5404 135614 5460
rect 135874 5404 135884 5460
rect 135940 5404 137340 5460
rect 137396 5404 137564 5460
rect 137620 5404 137630 5460
rect 14578 5292 14588 5348
rect 14644 5292 15820 5348
rect 15876 5292 15886 5348
rect 16034 5292 16044 5348
rect 16100 5292 18732 5348
rect 18788 5292 18798 5348
rect 40002 5292 40012 5348
rect 40068 5292 45948 5348
rect 46004 5292 46014 5348
rect 51202 5292 51212 5348
rect 51268 5292 53564 5348
rect 53620 5292 53630 5348
rect 62290 5292 62300 5348
rect 62356 5292 62748 5348
rect 62804 5292 66332 5348
rect 66388 5292 66398 5348
rect 71708 5236 71764 5404
rect 97412 5348 97468 5404
rect 132692 5348 132748 5404
rect 142044 5348 142100 5516
rect 158066 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158350 5516
rect 71922 5292 71932 5348
rect 71988 5292 75404 5348
rect 75460 5292 75470 5348
rect 75618 5292 75628 5348
rect 75684 5292 76972 5348
rect 77028 5292 78484 5348
rect 82674 5292 82684 5348
rect 82740 5292 83020 5348
rect 83076 5292 83086 5348
rect 84466 5292 84476 5348
rect 84532 5292 84542 5348
rect 89282 5292 89292 5348
rect 89348 5292 92092 5348
rect 92148 5292 92158 5348
rect 95340 5292 97468 5348
rect 101714 5292 101724 5348
rect 101780 5292 102060 5348
rect 102116 5292 102126 5348
rect 102386 5292 102396 5348
rect 102452 5292 103292 5348
rect 103348 5292 103358 5348
rect 105634 5292 105644 5348
rect 105700 5292 108556 5348
rect 108612 5292 108622 5348
rect 111458 5292 111468 5348
rect 111524 5292 112252 5348
rect 112308 5292 114940 5348
rect 114996 5292 115006 5348
rect 116050 5292 116060 5348
rect 116116 5292 117068 5348
rect 117124 5292 117516 5348
rect 117572 5292 117582 5348
rect 121650 5292 121660 5348
rect 121716 5292 122668 5348
rect 122724 5292 122734 5348
rect 123442 5292 123452 5348
rect 123508 5292 124460 5348
rect 124516 5292 132020 5348
rect 132672 5292 132748 5348
rect 132804 5292 133420 5348
rect 133476 5292 133486 5348
rect 135426 5292 135436 5348
rect 135492 5292 137676 5348
rect 137732 5292 137742 5348
rect 142044 5292 143948 5348
rect 144004 5292 144508 5348
rect 144564 5292 144574 5348
rect 147298 5292 147308 5348
rect 147364 5292 173180 5348
rect 173236 5292 173246 5348
rect 13682 5180 13692 5236
rect 13748 5180 14812 5236
rect 14868 5180 14878 5236
rect 15026 5180 15036 5236
rect 15092 5180 15102 5236
rect 19058 5180 19068 5236
rect 19124 5180 21644 5236
rect 21700 5180 21710 5236
rect 21858 5180 21868 5236
rect 21924 5180 23772 5236
rect 23828 5180 35644 5236
rect 35700 5180 37660 5236
rect 37716 5180 39228 5236
rect 39284 5180 39294 5236
rect 42578 5180 42588 5236
rect 42644 5180 45052 5236
rect 45108 5180 45118 5236
rect 49746 5180 49756 5236
rect 49812 5180 51436 5236
rect 51492 5180 51502 5236
rect 54562 5180 54572 5236
rect 54628 5180 57932 5236
rect 57988 5180 57998 5236
rect 58482 5180 58492 5236
rect 58548 5180 59500 5236
rect 59556 5180 59566 5236
rect 61628 5180 65660 5236
rect 65716 5180 67228 5236
rect 68226 5180 68236 5236
rect 68292 5180 69580 5236
rect 69636 5180 69646 5236
rect 71698 5180 71708 5236
rect 71764 5180 71774 5236
rect 7858 5068 7868 5124
rect 7924 5068 8652 5124
rect 8708 5068 8718 5124
rect 11666 5068 11676 5124
rect 11732 5068 12012 5124
rect 12068 5068 12078 5124
rect 12898 5068 12908 5124
rect 12964 5068 14252 5124
rect 14308 5068 14318 5124
rect 15036 5012 15092 5180
rect 61628 5124 61684 5180
rect 67172 5124 67228 5180
rect 73500 5124 73556 5292
rect 75282 5180 75292 5236
rect 75348 5180 76188 5236
rect 76244 5180 76254 5236
rect 78428 5124 78484 5292
rect 84476 5236 84532 5292
rect 95340 5236 95396 5292
rect 131964 5236 132020 5292
rect 78614 5180 78652 5236
rect 78708 5180 78718 5236
rect 81218 5180 81228 5236
rect 81284 5180 85484 5236
rect 85540 5180 85550 5236
rect 87938 5180 87948 5236
rect 88004 5180 88172 5236
rect 88228 5180 90412 5236
rect 90468 5180 90478 5236
rect 91298 5180 91308 5236
rect 91364 5180 92316 5236
rect 92372 5180 92382 5236
rect 94994 5180 95004 5236
rect 95060 5180 95340 5236
rect 95396 5180 95406 5236
rect 97122 5180 97132 5236
rect 97188 5180 98924 5236
rect 98980 5180 98990 5236
rect 99782 5180 99820 5236
rect 99876 5180 99886 5236
rect 101042 5180 101052 5236
rect 101108 5180 105420 5236
rect 105476 5180 105486 5236
rect 106306 5180 106316 5236
rect 106372 5180 113036 5236
rect 113092 5180 113102 5236
rect 119858 5180 119868 5236
rect 119924 5180 121716 5236
rect 121874 5180 121884 5236
rect 121940 5180 125020 5236
rect 125076 5180 125086 5236
rect 126018 5180 126028 5236
rect 126084 5180 127148 5236
rect 127204 5180 131740 5236
rect 131796 5180 131806 5236
rect 131964 5180 137788 5236
rect 137844 5180 137854 5236
rect 142258 5180 142268 5236
rect 142324 5180 147084 5236
rect 147140 5180 147644 5236
rect 147700 5180 147710 5236
rect 101052 5124 101108 5180
rect 121660 5124 121716 5180
rect 34850 5068 34860 5124
rect 34916 5068 35980 5124
rect 36036 5068 43260 5124
rect 43316 5068 43326 5124
rect 52546 5068 52556 5124
rect 52612 5068 53788 5124
rect 53844 5068 53854 5124
rect 57026 5068 57036 5124
rect 57092 5068 61684 5124
rect 61842 5068 61852 5124
rect 61908 5068 62860 5124
rect 62916 5068 62926 5124
rect 67172 5068 67676 5124
rect 67732 5068 67742 5124
rect 70214 5068 70252 5124
rect 70308 5068 70318 5124
rect 73490 5068 73500 5124
rect 73556 5068 73566 5124
rect 73826 5068 73836 5124
rect 73892 5068 75180 5124
rect 75236 5068 75246 5124
rect 75506 5068 75516 5124
rect 75572 5068 77644 5124
rect 77700 5068 77710 5124
rect 78428 5068 82292 5124
rect 88610 5068 88620 5124
rect 88676 5068 91084 5124
rect 91140 5068 91150 5124
rect 93212 5068 93772 5124
rect 93828 5068 93838 5124
rect 96310 5068 96348 5124
rect 96404 5068 96414 5124
rect 98802 5068 98812 5124
rect 98868 5068 101108 5124
rect 103730 5068 103740 5124
rect 103796 5068 105868 5124
rect 105924 5068 105934 5124
rect 109554 5068 109564 5124
rect 109620 5068 110236 5124
rect 110292 5068 114828 5124
rect 114884 5068 114894 5124
rect 115714 5068 115724 5124
rect 115780 5068 117404 5124
rect 117460 5068 117470 5124
rect 118514 5068 118524 5124
rect 118580 5068 118972 5124
rect 119028 5068 119038 5124
rect 119718 5068 119756 5124
rect 119812 5068 119822 5124
rect 120866 5068 120876 5124
rect 120932 5068 120942 5124
rect 121660 5068 122892 5124
rect 122948 5068 122958 5124
rect 123666 5068 123676 5124
rect 123732 5068 124908 5124
rect 124964 5068 124974 5124
rect 125346 5068 125356 5124
rect 125412 5068 127260 5124
rect 127316 5068 127326 5124
rect 127586 5068 127596 5124
rect 127652 5068 128156 5124
rect 128212 5068 128222 5124
rect 128482 5068 128492 5124
rect 128548 5068 131180 5124
rect 131236 5068 131246 5124
rect 133634 5068 133644 5124
rect 133700 5068 133980 5124
rect 134036 5068 134046 5124
rect 136098 5068 136108 5124
rect 136164 5068 136612 5124
rect 142034 5068 142044 5124
rect 142100 5068 144060 5124
rect 144116 5068 144126 5124
rect 82236 5012 82292 5068
rect 93212 5012 93268 5068
rect 118524 5012 118580 5068
rect 9874 4956 9884 5012
rect 9940 4956 14028 5012
rect 14084 4956 15092 5012
rect 31714 4956 31724 5012
rect 31780 4956 33908 5012
rect 35186 4956 35196 5012
rect 35252 4956 37996 5012
rect 38052 4956 38062 5012
rect 38210 4956 38220 5012
rect 38276 4956 38668 5012
rect 38724 4956 38734 5012
rect 40562 4956 40572 5012
rect 40628 4956 43036 5012
rect 43092 4956 43102 5012
rect 43922 4956 43932 5012
rect 43988 4956 48860 5012
rect 48916 4956 54012 5012
rect 54068 4956 54078 5012
rect 57138 4956 57148 5012
rect 57204 4956 60620 5012
rect 60676 4956 62356 5012
rect 62514 4956 62524 5012
rect 62580 4956 64316 5012
rect 64372 4956 64382 5012
rect 70466 4956 70476 5012
rect 70532 4956 71036 5012
rect 71092 4956 71102 5012
rect 71250 4956 71260 5012
rect 71316 4956 73612 5012
rect 73668 4956 73678 5012
rect 77074 4956 77084 5012
rect 77140 4956 77980 5012
rect 78036 4956 78046 5012
rect 78642 4956 78652 5012
rect 78708 4956 80220 5012
rect 80276 4956 81116 5012
rect 81172 4956 81182 5012
rect 82236 4956 83188 5012
rect 83458 4956 83468 5012
rect 83524 4956 84588 5012
rect 84644 4956 84654 5012
rect 89730 4956 89740 5012
rect 89796 4956 90972 5012
rect 91028 4956 91038 5012
rect 93202 4956 93212 5012
rect 93268 4956 93278 5012
rect 93650 4956 93660 5012
rect 93716 4956 94108 5012
rect 94164 4956 94174 5012
rect 96114 4956 96124 5012
rect 96180 4956 96796 5012
rect 96852 4956 96862 5012
rect 100370 4956 100380 5012
rect 100436 4956 102844 5012
rect 102900 4956 102910 5012
rect 104402 4956 104412 5012
rect 104468 4956 106540 5012
rect 106596 4956 106606 5012
rect 108322 4956 108332 5012
rect 108388 4956 108892 5012
rect 108948 4956 108958 5012
rect 111794 4956 111804 5012
rect 111860 4956 118580 5012
rect 120876 5012 120932 5068
rect 136556 5012 136612 5068
rect 120876 4956 121772 5012
rect 121828 4956 121838 5012
rect 122070 4956 122108 5012
rect 122164 4956 122174 5012
rect 124226 4956 124236 5012
rect 124292 4956 125132 5012
rect 125188 4956 125198 5012
rect 127698 4956 127708 5012
rect 127764 4956 130620 5012
rect 130676 4956 130686 5012
rect 133858 4956 133868 5012
rect 133924 4956 135100 5012
rect 135156 4956 135660 5012
rect 135716 4956 135726 5012
rect 136556 4956 136668 5012
rect 136724 4956 136734 5012
rect 137330 4956 137340 5012
rect 137396 4956 137900 5012
rect 137956 4956 137966 5012
rect 138338 4956 138348 5012
rect 138404 4956 138414 5012
rect 141250 4956 141260 5012
rect 141316 4956 145292 5012
rect 145348 4956 145516 5012
rect 145572 4956 146188 5012
rect 146244 4956 146748 5012
rect 146804 4956 146814 5012
rect 147746 4956 147756 5012
rect 147812 4956 147822 5012
rect 33852 4900 33908 4956
rect 62300 4900 62356 4956
rect 19170 4844 19180 4900
rect 19236 4844 32508 4900
rect 32564 4844 33516 4900
rect 33572 4844 33582 4900
rect 33842 4844 33852 4900
rect 33908 4844 35644 4900
rect 35700 4844 35710 4900
rect 36082 4844 36092 4900
rect 36148 4844 37548 4900
rect 37604 4844 37614 4900
rect 38994 4844 39004 4900
rect 39060 4844 40124 4900
rect 40180 4844 40190 4900
rect 43362 4844 43372 4900
rect 43428 4844 61404 4900
rect 61460 4844 61470 4900
rect 62300 4844 63196 4900
rect 63252 4844 64092 4900
rect 64148 4844 65772 4900
rect 65828 4844 65838 4900
rect 67442 4844 67452 4900
rect 67508 4844 67788 4900
rect 67844 4844 67854 4900
rect 68002 4844 68012 4900
rect 68068 4844 70364 4900
rect 70420 4844 70430 4900
rect 70802 4844 70812 4900
rect 70868 4844 72492 4900
rect 72548 4844 72558 4900
rect 76738 4844 76748 4900
rect 76804 4844 78092 4900
rect 78148 4844 78158 4900
rect 78418 4844 78428 4900
rect 78484 4844 79324 4900
rect 79380 4844 79390 4900
rect 80098 4844 80108 4900
rect 80164 4844 82964 4900
rect 36306 4732 36316 4788
rect 36372 4732 40572 4788
rect 40628 4732 40638 4788
rect 41570 4732 41580 4788
rect 41636 4732 44380 4788
rect 44436 4732 44446 4788
rect 64418 4732 64428 4788
rect 64484 4732 69132 4788
rect 69188 4732 69198 4788
rect 69346 4732 69356 4788
rect 69412 4732 70588 4788
rect 70644 4732 70654 4788
rect 76514 4732 76524 4788
rect 76580 4732 77308 4788
rect 77364 4732 78652 4788
rect 78708 4732 78718 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 81266 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81550 4732
rect 82908 4676 82964 4844
rect 83132 4788 83188 4956
rect 138348 4900 138404 4956
rect 147756 4900 147812 4956
rect 83318 4844 83356 4900
rect 83412 4844 83422 4900
rect 84018 4844 84028 4900
rect 84084 4844 84924 4900
rect 84980 4844 84990 4900
rect 85810 4844 85820 4900
rect 85876 4844 86604 4900
rect 86660 4844 89964 4900
rect 90020 4844 90188 4900
rect 90244 4844 90524 4900
rect 90580 4844 90590 4900
rect 91410 4844 91420 4900
rect 91476 4844 94668 4900
rect 94724 4844 94734 4900
rect 95330 4844 95340 4900
rect 95396 4844 96460 4900
rect 96516 4844 96526 4900
rect 97010 4844 97020 4900
rect 97076 4844 98812 4900
rect 98868 4844 98878 4900
rect 101266 4844 101276 4900
rect 101332 4844 102956 4900
rect 103012 4844 103022 4900
rect 103282 4844 103292 4900
rect 103348 4844 105980 4900
rect 106036 4844 106046 4900
rect 106204 4844 107548 4900
rect 107604 4844 107614 4900
rect 110562 4844 110572 4900
rect 110628 4844 113932 4900
rect 113988 4844 113998 4900
rect 115602 4844 115612 4900
rect 115668 4844 117516 4900
rect 117572 4844 119420 4900
rect 119476 4844 119486 4900
rect 121090 4844 121100 4900
rect 121156 4844 123340 4900
rect 123396 4844 123406 4900
rect 128146 4844 128156 4900
rect 128212 4844 129948 4900
rect 130004 4844 130844 4900
rect 130900 4844 130910 4900
rect 133746 4844 133756 4900
rect 133812 4844 138404 4900
rect 138786 4844 138796 4900
rect 138852 4844 139132 4900
rect 139188 4844 147812 4900
rect 149986 4844 149996 4900
rect 150052 4844 150668 4900
rect 150724 4844 150734 4900
rect 169250 4844 169260 4900
rect 169316 4844 169326 4900
rect 106204 4788 106260 4844
rect 83132 4732 84476 4788
rect 84532 4732 84542 4788
rect 85586 4732 85596 4788
rect 85652 4732 91308 4788
rect 91364 4732 91374 4788
rect 91634 4732 91644 4788
rect 91700 4732 104524 4788
rect 104580 4732 104590 4788
rect 105298 4732 105308 4788
rect 105364 4732 106260 4788
rect 107314 4732 107324 4788
rect 107380 4732 111804 4788
rect 111860 4732 111870 4788
rect 112578 4732 112588 4788
rect 112644 4732 113932 4788
rect 113988 4732 115948 4788
rect 116004 4732 116014 4788
rect 117618 4732 117628 4788
rect 117684 4732 121268 4788
rect 131058 4732 131068 4788
rect 131124 4732 133868 4788
rect 133924 4732 134652 4788
rect 134708 4732 135324 4788
rect 135380 4732 135390 4788
rect 135874 4732 135884 4788
rect 135940 4732 141596 4788
rect 141652 4732 141662 4788
rect 143714 4732 143724 4788
rect 143780 4732 145852 4788
rect 145908 4732 148652 4788
rect 148708 4732 148718 4788
rect 111986 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112270 4732
rect 121212 4676 121268 4732
rect 142706 4676 142716 4732
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142980 4676 142990 4732
rect 51986 4620 51996 4676
rect 52052 4620 57708 4676
rect 57764 4620 57774 4676
rect 62262 4620 62300 4676
rect 62356 4620 65212 4676
rect 65268 4620 66444 4676
rect 66500 4620 66510 4676
rect 66658 4620 66668 4676
rect 66724 4620 68124 4676
rect 68180 4620 68190 4676
rect 68898 4620 68908 4676
rect 68964 4620 76356 4676
rect 77382 4620 77420 4676
rect 77476 4620 77486 4676
rect 82908 4620 91308 4676
rect 91364 4620 91374 4676
rect 91532 4620 98476 4676
rect 98532 4620 98542 4676
rect 100258 4620 100268 4676
rect 100324 4620 109900 4676
rect 109956 4620 110460 4676
rect 110516 4620 110526 4676
rect 113362 4620 113372 4676
rect 113428 4620 115724 4676
rect 115780 4620 120932 4676
rect 121202 4620 121212 4676
rect 121268 4620 121436 4676
rect 121492 4620 121502 4676
rect 123554 4620 123564 4676
rect 123620 4620 123900 4676
rect 123956 4620 123966 4676
rect 129266 4620 129276 4676
rect 129332 4620 129724 4676
rect 129780 4620 130844 4676
rect 130900 4620 130910 4676
rect 133074 4620 133084 4676
rect 133140 4620 133756 4676
rect 133812 4620 133822 4676
rect 136770 4620 136780 4676
rect 136836 4620 139692 4676
rect 139748 4620 139758 4676
rect 140914 4620 140924 4676
rect 140980 4620 142156 4676
rect 142212 4620 142222 4676
rect 143266 4620 143276 4676
rect 143332 4620 145180 4676
rect 145236 4620 145246 4676
rect 10434 4508 10444 4564
rect 10500 4508 31948 4564
rect 33506 4508 33516 4564
rect 33572 4508 39452 4564
rect 39508 4508 39518 4564
rect 40786 4508 40796 4564
rect 40852 4508 58940 4564
rect 58996 4508 59006 4564
rect 59500 4508 60956 4564
rect 61012 4508 61022 4564
rect 61842 4508 61852 4564
rect 61908 4508 70756 4564
rect 71362 4508 71372 4564
rect 71428 4508 73612 4564
rect 73668 4508 73678 4564
rect 17154 4396 17164 4452
rect 17220 4396 18396 4452
rect 18452 4396 18462 4452
rect 23426 4396 23436 4452
rect 23492 4396 27580 4452
rect 27636 4396 28588 4452
rect 28644 4396 28654 4452
rect 31892 4340 31948 4508
rect 59500 4452 59556 4508
rect 40674 4396 40684 4452
rect 40740 4396 42364 4452
rect 42420 4396 42430 4452
rect 43250 4396 43260 4452
rect 43316 4396 59556 4452
rect 59714 4396 59724 4452
rect 59780 4396 60508 4452
rect 60564 4396 60574 4452
rect 62066 4396 62076 4452
rect 62132 4396 64428 4452
rect 64484 4396 64494 4452
rect 64642 4396 64652 4452
rect 64708 4396 64718 4452
rect 67106 4396 67116 4452
rect 67172 4396 67900 4452
rect 67956 4396 67966 4452
rect 68310 4396 68348 4452
rect 68404 4396 68414 4452
rect 69122 4396 69132 4452
rect 69188 4396 70644 4452
rect 64652 4340 64708 4396
rect 22866 4284 22876 4340
rect 22932 4284 23324 4340
rect 23380 4284 25340 4340
rect 25396 4284 25406 4340
rect 31892 4284 32844 4340
rect 32900 4284 40348 4340
rect 40404 4284 40414 4340
rect 40786 4284 40796 4340
rect 40852 4284 42252 4340
rect 42308 4284 42318 4340
rect 42578 4284 42588 4340
rect 42644 4284 43148 4340
rect 43204 4284 43214 4340
rect 43652 4284 45388 4340
rect 45444 4284 48412 4340
rect 48468 4284 51996 4340
rect 52052 4284 52062 4340
rect 57474 4284 57484 4340
rect 57540 4284 62524 4340
rect 62580 4284 62590 4340
rect 64652 4284 69356 4340
rect 69412 4284 69422 4340
rect 43652 4228 43708 4284
rect 70588 4228 70644 4396
rect 70700 4340 70756 4508
rect 76300 4452 76356 4620
rect 76514 4508 76524 4564
rect 76580 4508 82236 4564
rect 82292 4508 83356 4564
rect 83412 4508 83422 4564
rect 83794 4508 83804 4564
rect 83860 4508 85148 4564
rect 85204 4508 85214 4564
rect 88386 4508 88396 4564
rect 88452 4508 88844 4564
rect 88900 4508 90076 4564
rect 90132 4508 90142 4564
rect 91532 4452 91588 4620
rect 120876 4564 120932 4620
rect 92418 4508 92428 4564
rect 92484 4508 93324 4564
rect 93380 4508 93390 4564
rect 95106 4508 95116 4564
rect 95172 4508 97020 4564
rect 97076 4508 97086 4564
rect 102162 4508 102172 4564
rect 102228 4508 105308 4564
rect 105364 4508 105374 4564
rect 106418 4508 106428 4564
rect 106484 4508 113092 4564
rect 113222 4508 113260 4564
rect 113316 4508 113326 4564
rect 113698 4508 113708 4564
rect 113764 4508 116060 4564
rect 116116 4508 116126 4564
rect 117282 4508 117292 4564
rect 117348 4508 117404 4564
rect 117460 4508 117470 4564
rect 118188 4508 120484 4564
rect 120866 4508 120876 4564
rect 120932 4508 121324 4564
rect 121380 4508 121390 4564
rect 121650 4508 121660 4564
rect 121716 4508 126812 4564
rect 126868 4508 126878 4564
rect 127698 4508 127708 4564
rect 127764 4508 127932 4564
rect 127988 4508 127998 4564
rect 129052 4508 131628 4564
rect 131684 4508 131694 4564
rect 135622 4508 135660 4564
rect 135716 4508 135726 4564
rect 135874 4508 135884 4564
rect 135940 4508 135978 4564
rect 138562 4508 138572 4564
rect 138628 4508 141708 4564
rect 141764 4508 141774 4564
rect 143042 4508 143052 4564
rect 143108 4508 144060 4564
rect 144116 4508 144126 4564
rect 147634 4508 147644 4564
rect 147700 4508 148764 4564
rect 148820 4508 149100 4564
rect 149156 4508 149166 4564
rect 70914 4396 70924 4452
rect 70980 4396 71820 4452
rect 71876 4396 71886 4452
rect 72594 4396 72604 4452
rect 72660 4396 74060 4452
rect 74116 4396 74126 4452
rect 76300 4396 78204 4452
rect 78260 4396 78270 4452
rect 82338 4396 82348 4452
rect 82404 4396 84252 4452
rect 84308 4396 84318 4452
rect 84802 4396 84812 4452
rect 84868 4396 91588 4452
rect 92978 4396 92988 4452
rect 93044 4396 96348 4452
rect 96404 4396 96414 4452
rect 96786 4396 96796 4452
rect 96852 4396 97356 4452
rect 97412 4396 101500 4452
rect 101556 4396 101566 4452
rect 103282 4396 103292 4452
rect 103348 4396 104188 4452
rect 104244 4396 104254 4452
rect 104738 4396 104748 4452
rect 104804 4396 111356 4452
rect 111412 4396 111422 4452
rect 113036 4340 113092 4508
rect 114594 4396 114604 4452
rect 114660 4396 116172 4452
rect 116228 4396 116238 4452
rect 70700 4284 72380 4340
rect 72436 4284 72940 4340
rect 72996 4284 73006 4340
rect 74386 4284 74396 4340
rect 74452 4284 74956 4340
rect 75012 4284 75022 4340
rect 82898 4284 82908 4340
rect 82964 4284 83804 4340
rect 83860 4284 83870 4340
rect 85558 4284 85596 4340
rect 85652 4284 85662 4340
rect 89394 4284 89404 4340
rect 89460 4284 92540 4340
rect 92596 4284 92764 4340
rect 92820 4284 92830 4340
rect 102134 4284 102172 4340
rect 102228 4284 102238 4340
rect 104178 4284 104188 4340
rect 104244 4284 105420 4340
rect 105476 4284 105486 4340
rect 105970 4284 105980 4340
rect 106036 4284 108108 4340
rect 108164 4284 111468 4340
rect 111524 4284 111534 4340
rect 113036 4284 117964 4340
rect 118020 4284 118030 4340
rect 85596 4228 85652 4284
rect 118188 4228 118244 4508
rect 120428 4452 120484 4508
rect 129052 4452 129108 4508
rect 169260 4452 169316 4844
rect 173426 4676 173436 4732
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173700 4676 173710 4732
rect 119410 4396 119420 4452
rect 119476 4396 120204 4452
rect 120260 4396 120270 4452
rect 120428 4396 121548 4452
rect 121604 4396 121614 4452
rect 125794 4396 125804 4452
rect 125860 4396 129052 4452
rect 129108 4396 129118 4452
rect 131058 4396 131068 4452
rect 131124 4396 136108 4452
rect 136164 4396 136174 4452
rect 148082 4396 148092 4452
rect 148148 4396 149660 4452
rect 149716 4396 149726 4452
rect 150780 4396 157388 4452
rect 157444 4396 157454 4452
rect 169250 4396 169260 4452
rect 169316 4396 169326 4452
rect 150780 4340 150836 4396
rect 118850 4284 118860 4340
rect 118916 4284 119868 4340
rect 119924 4284 119934 4340
rect 121202 4284 121212 4340
rect 121268 4284 121324 4340
rect 121380 4284 121390 4340
rect 122322 4284 122332 4340
rect 122388 4284 126252 4340
rect 126308 4284 126318 4340
rect 128034 4284 128044 4340
rect 128100 4284 128716 4340
rect 128772 4284 128782 4340
rect 132402 4284 132412 4340
rect 132468 4284 134428 4340
rect 134484 4284 134494 4340
rect 138674 4284 138684 4340
rect 138740 4284 140252 4340
rect 140308 4284 140588 4340
rect 140644 4284 140654 4340
rect 141810 4284 141820 4340
rect 141876 4284 145068 4340
rect 145124 4284 145134 4340
rect 147298 4284 147308 4340
rect 147364 4284 147374 4340
rect 149090 4284 149100 4340
rect 149156 4284 149772 4340
rect 149828 4284 150836 4340
rect 150994 4284 151004 4340
rect 151060 4284 151452 4340
rect 151508 4284 151518 4340
rect 161074 4284 161084 4340
rect 161140 4284 161532 4340
rect 161588 4284 161598 4340
rect 147308 4228 147364 4284
rect 9090 4172 9100 4228
rect 9156 4172 9884 4228
rect 9940 4172 9950 4228
rect 16146 4172 16156 4228
rect 16212 4172 17836 4228
rect 17892 4172 28588 4228
rect 28644 4172 29148 4228
rect 29204 4172 38668 4228
rect 38724 4172 41692 4228
rect 41748 4172 43708 4228
rect 44370 4172 44380 4228
rect 44436 4172 50876 4228
rect 50932 4172 50942 4228
rect 54674 4172 54684 4228
rect 54740 4172 55580 4228
rect 55636 4172 55646 4228
rect 64866 4172 64876 4228
rect 64932 4172 66108 4228
rect 66164 4172 66174 4228
rect 69234 4172 69244 4228
rect 69300 4172 70028 4228
rect 70084 4172 70094 4228
rect 70588 4172 76300 4228
rect 76356 4172 76366 4228
rect 77970 4172 77980 4228
rect 78036 4172 85652 4228
rect 90962 4172 90972 4228
rect 91028 4172 92204 4228
rect 92260 4172 93772 4228
rect 93828 4172 93838 4228
rect 97794 4172 97804 4228
rect 97860 4172 98700 4228
rect 98756 4172 98766 4228
rect 106194 4172 106204 4228
rect 106260 4172 107100 4228
rect 107156 4172 107166 4228
rect 107538 4172 107548 4228
rect 107604 4172 108444 4228
rect 108500 4172 108510 4228
rect 109554 4172 109564 4228
rect 109620 4172 110236 4228
rect 110292 4172 110302 4228
rect 114454 4172 114492 4228
rect 114548 4172 114558 4228
rect 115154 4172 115164 4228
rect 115220 4172 115500 4228
rect 115556 4172 118244 4228
rect 118626 4172 118636 4228
rect 118692 4172 120988 4228
rect 122210 4172 122220 4228
rect 122276 4172 124796 4228
rect 124852 4172 125692 4228
rect 125748 4172 125758 4228
rect 133830 4172 133868 4228
rect 133924 4172 133934 4228
rect 134642 4172 134652 4228
rect 134708 4172 137116 4228
rect 137172 4172 139468 4228
rect 139524 4172 139692 4228
rect 139748 4172 139758 4228
rect 142258 4172 142268 4228
rect 142324 4172 143052 4228
rect 143108 4172 143118 4228
rect 143490 4172 143500 4228
rect 143556 4172 143724 4228
rect 143780 4172 143790 4228
rect 147308 4172 151676 4228
rect 151732 4172 151742 4228
rect 6850 4060 6860 4116
rect 6916 4060 8540 4116
rect 8596 4060 35868 4116
rect 35924 4060 35934 4116
rect 39890 4060 39900 4116
rect 39956 4060 40796 4116
rect 40852 4060 40862 4116
rect 63634 4060 63644 4116
rect 63700 4060 74620 4116
rect 74676 4060 74686 4116
rect 89170 4060 89180 4116
rect 89236 4060 91756 4116
rect 91812 4060 91822 4116
rect 96898 4060 96908 4116
rect 96964 4060 98924 4116
rect 98980 4060 98990 4116
rect 109442 4060 109452 4116
rect 109508 4060 116956 4116
rect 117012 4060 117022 4116
rect 120932 4004 120988 4172
rect 121538 4060 121548 4116
rect 121604 4060 122668 4116
rect 122724 4060 122734 4116
rect 123554 4060 123564 4116
rect 123620 4060 124124 4116
rect 124180 4060 124190 4116
rect 125122 4060 125132 4116
rect 125188 4060 129164 4116
rect 129220 4060 129230 4116
rect 138562 4060 138572 4116
rect 138628 4060 140476 4116
rect 140532 4060 148652 4116
rect 148708 4060 148718 4116
rect 15810 3948 15820 4004
rect 15876 3948 17724 4004
rect 17780 3948 17790 4004
rect 39666 3948 39676 4004
rect 39732 3948 64764 4004
rect 64820 3948 64830 4004
rect 76290 3948 76300 4004
rect 76356 3948 77252 4004
rect 80434 3948 80444 4004
rect 80500 3948 91980 4004
rect 92036 3948 92046 4004
rect 120932 3948 123228 4004
rect 123284 3948 123294 4004
rect 128594 3948 128604 4004
rect 128660 3948 132188 4004
rect 132244 3948 132254 4004
rect 134306 3948 134316 4004
rect 134372 3948 137340 4004
rect 137396 3948 137564 4004
rect 137620 3948 137630 4004
rect 137778 3948 137788 4004
rect 137844 3948 141148 4004
rect 141204 3948 141214 4004
rect 144274 3948 144284 4004
rect 144340 3948 146300 4004
rect 146356 3948 146366 4004
rect 149762 3948 149772 4004
rect 149828 3948 151116 4004
rect 151172 3948 151182 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 77196 3892 77252 3948
rect 96626 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96910 3948
rect 127346 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127630 3948
rect 158066 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158350 3948
rect 73892 3836 74844 3892
rect 74900 3836 76972 3892
rect 77028 3836 77038 3892
rect 77196 3836 85708 3892
rect 108434 3836 108444 3892
rect 108500 3836 116396 3892
rect 116452 3836 116462 3892
rect 119634 3836 119644 3892
rect 119700 3836 121436 3892
rect 121492 3836 121502 3892
rect 121762 3836 121772 3892
rect 121828 3836 123676 3892
rect 123732 3836 123742 3892
rect 124114 3836 124124 3892
rect 124180 3836 126140 3892
rect 126196 3836 126700 3892
rect 126756 3836 126766 3892
rect 128034 3836 128044 3892
rect 128100 3836 129836 3892
rect 129892 3836 129902 3892
rect 130274 3836 130284 3892
rect 130340 3836 132636 3892
rect 132692 3836 132702 3892
rect 136322 3836 136332 3892
rect 136388 3836 138908 3892
rect 138964 3836 138974 3892
rect 148194 3836 148204 3892
rect 148260 3836 150556 3892
rect 150612 3836 150622 3892
rect 150892 3836 156492 3892
rect 156548 3836 156558 3892
rect 73892 3780 73948 3836
rect 85652 3780 85708 3836
rect 150892 3780 150948 3836
rect 11442 3724 11452 3780
rect 11508 3724 20188 3780
rect 25442 3724 25452 3780
rect 25508 3724 27132 3780
rect 27188 3724 27198 3780
rect 29474 3724 29484 3780
rect 29540 3724 30044 3780
rect 30100 3724 32284 3780
rect 32340 3724 32350 3780
rect 41020 3724 42588 3780
rect 42644 3724 42654 3780
rect 46162 3724 46172 3780
rect 46228 3724 46238 3780
rect 63522 3724 63532 3780
rect 63588 3724 66108 3780
rect 66164 3724 66174 3780
rect 67172 3724 73948 3780
rect 75954 3724 75964 3780
rect 76020 3724 76860 3780
rect 76916 3724 76926 3780
rect 79314 3724 79324 3780
rect 79380 3724 79996 3780
rect 80052 3724 80062 3780
rect 85652 3724 92652 3780
rect 92708 3724 92718 3780
rect 94434 3724 94444 3780
rect 94500 3724 95340 3780
rect 95396 3724 95406 3780
rect 102386 3724 102396 3780
rect 102452 3724 110796 3780
rect 110852 3724 110862 3780
rect 120194 3724 120204 3780
rect 120260 3724 121548 3780
rect 121604 3724 121614 3780
rect 127586 3724 127596 3780
rect 127652 3724 130060 3780
rect 130116 3724 130126 3780
rect 130508 3724 132972 3780
rect 133028 3724 133420 3780
rect 133476 3724 133486 3780
rect 133746 3724 133756 3780
rect 133812 3724 136220 3780
rect 136276 3724 137116 3780
rect 137172 3724 137182 3780
rect 137330 3724 137340 3780
rect 137396 3724 138012 3780
rect 138068 3724 138078 3780
rect 138460 3724 139020 3780
rect 139076 3724 139086 3780
rect 140466 3724 140476 3780
rect 140532 3724 143276 3780
rect 143332 3724 143836 3780
rect 143892 3724 143902 3780
rect 145170 3724 145180 3780
rect 145236 3724 145628 3780
rect 145684 3724 145694 3780
rect 148866 3724 148876 3780
rect 148932 3724 149996 3780
rect 150052 3724 150062 3780
rect 150220 3724 150948 3780
rect 151106 3724 151116 3780
rect 151172 3724 152012 3780
rect 152068 3724 152078 3780
rect 20132 3668 20188 3724
rect 41020 3668 41076 3724
rect 12114 3612 12124 3668
rect 12180 3612 13804 3668
rect 13860 3612 19292 3668
rect 19348 3612 19358 3668
rect 20132 3612 41076 3668
rect 41234 3612 41244 3668
rect 41300 3612 41804 3668
rect 41860 3612 41870 3668
rect 46172 3556 46228 3724
rect 67172 3668 67228 3724
rect 130508 3668 130564 3724
rect 64754 3612 64764 3668
rect 64820 3612 67228 3668
rect 73602 3612 73612 3668
rect 73668 3612 77084 3668
rect 77140 3612 77532 3668
rect 77588 3612 77598 3668
rect 94770 3612 94780 3668
rect 94836 3612 97468 3668
rect 104738 3612 104748 3668
rect 104804 3612 109116 3668
rect 109172 3612 109182 3668
rect 112914 3612 112924 3668
rect 112980 3612 114044 3668
rect 114100 3612 114110 3668
rect 116274 3612 116284 3668
rect 116340 3612 117964 3668
rect 118020 3612 118030 3668
rect 120754 3612 120764 3668
rect 120820 3612 121604 3668
rect 121874 3612 121884 3668
rect 121940 3612 125356 3668
rect 125412 3612 125422 3668
rect 125794 3612 125804 3668
rect 125860 3612 128492 3668
rect 128548 3612 128558 3668
rect 129154 3612 129164 3668
rect 129220 3612 130564 3668
rect 130620 3612 131292 3668
rect 131348 3612 131516 3668
rect 131572 3612 131582 3668
rect 132178 3612 132188 3668
rect 132244 3612 135212 3668
rect 135268 3612 135436 3668
rect 135492 3612 135502 3668
rect 97412 3556 97468 3612
rect 121548 3556 121604 3612
rect 130620 3556 130676 3612
rect 138460 3556 138516 3724
rect 14242 3500 14252 3556
rect 14308 3500 14700 3556
rect 14756 3500 16604 3556
rect 16660 3500 16670 3556
rect 20626 3500 20636 3556
rect 20692 3500 21980 3556
rect 22036 3500 22428 3556
rect 22484 3500 22494 3556
rect 24098 3500 24108 3556
rect 24164 3500 24556 3556
rect 24612 3500 27244 3556
rect 27300 3500 27310 3556
rect 28242 3500 28252 3556
rect 28308 3500 29260 3556
rect 29316 3500 30604 3556
rect 30660 3500 30670 3556
rect 45490 3500 45500 3556
rect 45556 3500 46844 3556
rect 46900 3500 46910 3556
rect 65538 3500 65548 3556
rect 65604 3500 68460 3556
rect 68516 3500 68526 3556
rect 88050 3500 88060 3556
rect 88116 3500 89628 3556
rect 89684 3500 89694 3556
rect 92754 3500 92764 3556
rect 92820 3500 94668 3556
rect 94724 3500 94734 3556
rect 97412 3500 98476 3556
rect 98532 3500 107548 3556
rect 107604 3500 107614 3556
rect 112354 3500 112364 3556
rect 112420 3500 113372 3556
rect 113428 3500 113438 3556
rect 121174 3500 121212 3556
rect 121268 3500 121278 3556
rect 121548 3500 124348 3556
rect 124404 3500 124414 3556
rect 125234 3500 125244 3556
rect 125300 3500 127036 3556
rect 127092 3500 127260 3556
rect 127316 3500 127326 3556
rect 127474 3500 127484 3556
rect 127540 3500 130676 3556
rect 130834 3500 130844 3556
rect 130900 3500 133644 3556
rect 133700 3500 134204 3556
rect 134260 3500 134270 3556
rect 135314 3500 135324 3556
rect 135380 3500 138516 3556
rect 138684 3612 139972 3668
rect 142594 3612 142604 3668
rect 142660 3612 144732 3668
rect 144788 3612 144956 3668
rect 145012 3612 145022 3668
rect 146066 3612 146076 3668
rect 146132 3612 147532 3668
rect 147588 3612 148092 3668
rect 148148 3612 148158 3668
rect 149314 3612 149324 3668
rect 149380 3612 149772 3668
rect 149828 3612 149838 3668
rect 138684 3444 138740 3612
rect 139916 3556 139972 3612
rect 150220 3556 150276 3724
rect 151900 3612 152796 3668
rect 152852 3612 152862 3668
rect 154354 3612 154364 3668
rect 154420 3612 155372 3668
rect 155428 3612 155820 3668
rect 155876 3612 155886 3668
rect 167794 3612 167804 3668
rect 167860 3612 169484 3668
rect 169540 3612 169550 3668
rect 151900 3556 151956 3612
rect 139906 3500 139916 3556
rect 139972 3500 140252 3556
rect 140308 3500 140318 3556
rect 142146 3500 142156 3556
rect 142212 3500 143612 3556
rect 143668 3500 144172 3556
rect 144228 3500 144238 3556
rect 145394 3500 145404 3556
rect 145460 3500 147196 3556
rect 147252 3500 147262 3556
rect 148978 3500 148988 3556
rect 149044 3500 150276 3556
rect 150434 3500 150444 3556
rect 150500 3500 151900 3556
rect 151956 3500 151966 3556
rect 152674 3500 152684 3556
rect 152740 3500 153692 3556
rect 153748 3500 154028 3556
rect 154084 3500 154094 3556
rect 155474 3500 155484 3556
rect 155540 3500 156716 3556
rect 156772 3500 156782 3556
rect 157714 3500 157724 3556
rect 157780 3500 158508 3556
rect 158564 3500 158956 3556
rect 159012 3500 159022 3556
rect 159394 3500 159404 3556
rect 159460 3500 160636 3556
rect 160692 3500 160702 3556
rect 162754 3500 162764 3556
rect 162820 3500 163660 3556
rect 163716 3500 164108 3556
rect 164164 3500 164174 3556
rect 164434 3500 164444 3556
rect 164500 3500 165452 3556
rect 165508 3500 165788 3556
rect 165844 3500 165854 3556
rect 166114 3500 166124 3556
rect 166180 3500 167132 3556
rect 167188 3500 167580 3556
rect 167636 3500 167646 3556
rect 169586 3500 169596 3556
rect 169652 3500 170716 3556
rect 170772 3500 170782 3556
rect 171154 3500 171164 3556
rect 171220 3500 172396 3556
rect 172452 3500 172462 3556
rect 5842 3388 5852 3444
rect 5908 3388 6524 3444
rect 6580 3388 6590 3444
rect 11218 3388 11228 3444
rect 11284 3388 11788 3444
rect 11844 3388 12124 3444
rect 12180 3388 12190 3444
rect 14802 3388 14812 3444
rect 14868 3388 16044 3444
rect 16100 3388 16110 3444
rect 17154 3388 17164 3444
rect 17220 3388 17836 3444
rect 17892 3388 17902 3444
rect 19730 3388 19740 3444
rect 19796 3388 21084 3444
rect 21140 3388 21150 3444
rect 23650 3388 23660 3444
rect 23716 3388 26124 3444
rect 26180 3388 26190 3444
rect 27458 3388 27468 3444
rect 27524 3388 28140 3444
rect 28196 3388 30492 3444
rect 30548 3388 30940 3444
rect 30996 3388 31006 3444
rect 31490 3388 31500 3444
rect 31556 3388 32060 3444
rect 32116 3388 32126 3444
rect 32834 3388 32844 3444
rect 32900 3388 33516 3444
rect 33572 3388 33582 3444
rect 35410 3388 35420 3444
rect 35476 3388 36204 3444
rect 36260 3388 36270 3444
rect 45378 3388 45388 3444
rect 45444 3388 46340 3444
rect 47730 3388 47740 3444
rect 47796 3388 49644 3444
rect 49700 3388 49710 3444
rect 55010 3388 55020 3444
rect 55076 3388 56364 3444
rect 56420 3388 56430 3444
rect 57138 3388 57148 3444
rect 57204 3388 58044 3444
rect 58100 3388 58110 3444
rect 58930 3388 58940 3444
rect 58996 3388 59724 3444
rect 59780 3388 59790 3444
rect 65874 3388 65884 3444
rect 65940 3388 67004 3444
rect 67060 3388 67070 3444
rect 67554 3388 67564 3444
rect 67620 3388 69356 3444
rect 69412 3388 69422 3444
rect 74386 3388 74396 3444
rect 74452 3388 75180 3444
rect 75236 3388 75246 3444
rect 77634 3388 77644 3444
rect 77700 3388 78764 3444
rect 78820 3388 78830 3444
rect 84354 3388 84364 3444
rect 84420 3388 85148 3444
rect 85204 3388 85214 3444
rect 89394 3388 89404 3444
rect 89460 3388 90524 3444
rect 90580 3388 90590 3444
rect 91074 3388 91084 3444
rect 91140 3388 92876 3444
rect 92932 3388 92942 3444
rect 96114 3388 96124 3444
rect 96180 3388 97244 3444
rect 97300 3388 97310 3444
rect 99474 3388 99484 3444
rect 99540 3388 100716 3444
rect 100772 3388 100782 3444
rect 101154 3388 101164 3444
rect 101220 3388 101948 3444
rect 102004 3388 102014 3444
rect 102844 3388 104076 3444
rect 104132 3388 104142 3444
rect 104514 3388 104524 3444
rect 104580 3388 106428 3444
rect 106484 3388 106494 3444
rect 107874 3388 107884 3444
rect 107940 3388 109004 3444
rect 109060 3388 109070 3444
rect 111234 3388 111244 3444
rect 111300 3388 111916 3444
rect 111972 3388 111982 3444
rect 114594 3388 114604 3444
rect 114660 3388 116396 3444
rect 116452 3388 116462 3444
rect 117954 3388 117964 3444
rect 118020 3388 120316 3444
rect 120372 3388 120382 3444
rect 120978 3388 120988 3444
rect 121044 3388 121772 3444
rect 121828 3388 121838 3444
rect 123554 3388 123564 3444
rect 123620 3388 126364 3444
rect 126420 3388 126430 3444
rect 126914 3388 126924 3444
rect 126980 3388 128940 3444
rect 128996 3388 129006 3444
rect 130162 3388 130172 3444
rect 130228 3388 130956 3444
rect 131012 3388 131022 3444
rect 132514 3388 132524 3444
rect 132580 3388 136332 3444
rect 136388 3388 136398 3444
rect 136994 3388 137004 3444
rect 137060 3388 138740 3444
rect 139122 3388 139132 3444
rect 139188 3388 142044 3444
rect 142100 3388 142110 3444
rect 143714 3388 143724 3444
rect 143780 3388 145292 3444
rect 145348 3388 145964 3444
rect 146020 3388 146030 3444
rect 147074 3388 147084 3444
rect 147140 3388 149884 3444
rect 149940 3388 149950 3444
rect 152114 3388 152124 3444
rect 152180 3388 152460 3444
rect 152516 3388 152908 3444
rect 152964 3388 152974 3444
rect 153906 3388 153916 3444
rect 153972 3388 154588 3444
rect 154644 3388 155036 3444
rect 155092 3388 155102 3444
rect 156594 3388 156604 3444
rect 156660 3388 157164 3444
rect 157220 3388 157230 3444
rect 158834 3388 158844 3444
rect 158900 3388 159292 3444
rect 159348 3388 159852 3444
rect 159908 3388 159918 3444
rect 160514 3388 160524 3444
rect 160580 3388 161644 3444
rect 161700 3388 161710 3444
rect 162194 3388 162204 3444
rect 162260 3388 162876 3444
rect 162932 3388 162942 3444
rect 163874 3388 163884 3444
rect 163940 3388 164668 3444
rect 164724 3388 164734 3444
rect 165666 3388 165676 3444
rect 165732 3388 166348 3444
rect 166404 3388 166796 3444
rect 166852 3388 166862 3444
rect 167234 3388 167244 3444
rect 167300 3388 168140 3444
rect 168196 3388 168588 3444
rect 168644 3388 168654 3444
rect 170594 3388 170604 3444
rect 170660 3388 171388 3444
rect 171444 3388 171612 3444
rect 171668 3388 171678 3444
rect 172274 3388 172284 3444
rect 172340 3388 173404 3444
rect 173460 3388 173470 3444
rect 46284 3332 46340 3388
rect 102844 3332 102900 3388
rect 14578 3276 14588 3332
rect 14644 3276 41356 3332
rect 41412 3276 41422 3332
rect 46274 3276 46284 3332
rect 46340 3276 46350 3332
rect 58370 3276 58380 3332
rect 58436 3276 61516 3332
rect 61572 3276 61582 3332
rect 96226 3276 96236 3332
rect 96292 3276 98140 3332
rect 98196 3276 100044 3332
rect 100100 3276 101836 3332
rect 101892 3276 101902 3332
rect 102834 3276 102844 3332
rect 102900 3276 102910 3332
rect 104626 3276 104636 3332
rect 104692 3276 118076 3332
rect 118132 3276 118142 3332
rect 119634 3276 119644 3332
rect 119700 3276 122444 3332
rect 122500 3276 122510 3332
rect 124198 3276 124236 3332
rect 124292 3276 124302 3332
rect 125570 3276 125580 3332
rect 125636 3276 126028 3332
rect 126084 3276 126094 3332
rect 128118 3276 128156 3332
rect 128212 3276 128222 3332
rect 131842 3276 131852 3332
rect 131908 3276 136892 3332
rect 136948 3276 136958 3332
rect 137732 3276 140364 3332
rect 140420 3276 140430 3332
rect 141484 3276 142940 3332
rect 142996 3276 143006 3332
rect 143938 3276 143948 3332
rect 144004 3276 146860 3332
rect 146916 3276 146926 3332
rect 147970 3276 147980 3332
rect 148036 3276 154700 3332
rect 154756 3276 154766 3332
rect 159170 3276 159180 3332
rect 159236 3276 165228 3332
rect 165284 3276 165294 3332
rect 173954 3276 173964 3332
rect 174020 3276 174972 3332
rect 175028 3276 175038 3332
rect 137732 3220 137788 3276
rect 141484 3220 141540 3276
rect 94098 3164 94108 3220
rect 94164 3164 106876 3220
rect 106932 3164 106942 3220
rect 122546 3164 122556 3220
rect 122612 3164 125132 3220
rect 125188 3164 125198 3220
rect 127810 3164 127820 3220
rect 127876 3164 129500 3220
rect 129556 3164 130060 3220
rect 130116 3164 130126 3220
rect 131954 3164 131964 3220
rect 132020 3164 137788 3220
rect 140130 3164 140140 3220
rect 140196 3164 141540 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 81266 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81550 3164
rect 111986 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112270 3164
rect 142706 3108 142716 3164
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142980 3108 142990 3164
rect 173426 3108 173436 3164
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173700 3108 173710 3164
rect 120082 3052 120092 3108
rect 120148 3052 127036 3108
rect 127092 3052 134092 3108
rect 134148 3052 134158 3108
rect 135762 3052 135772 3108
rect 135828 3052 139916 3108
rect 139972 3052 139982 3108
rect 39106 2940 39116 2996
rect 39172 2940 117292 2996
rect 117348 2940 117358 2996
rect 124898 2940 124908 2996
rect 124964 2940 150780 2996
rect 150836 2940 150846 2996
rect 52098 2828 52108 2884
rect 52164 2828 119196 2884
rect 119252 2828 119262 2884
rect 126130 2828 126140 2884
rect 126196 2828 139244 2884
rect 139300 2828 139310 2884
rect 141026 2828 141036 2884
rect 141092 2828 143836 2884
rect 143892 2828 143902 2884
rect 18162 2716 18172 2772
rect 18228 2716 57036 2772
rect 57092 2716 57102 2772
rect 93314 2716 93324 2772
rect 93380 2716 112700 2772
rect 112756 2716 112766 2772
rect 130498 2716 130508 2772
rect 130564 2716 168252 2772
rect 168308 2716 168318 2772
rect 11666 2604 11676 2660
rect 11732 2604 58380 2660
rect 58436 2604 58446 2660
rect 74610 2604 74620 2660
rect 74676 2604 132972 2660
rect 133028 2604 133038 2660
rect 136658 2604 136668 2660
rect 136724 2604 147308 2660
rect 147364 2604 147374 2660
rect 74722 2492 74732 2548
rect 74788 2492 131180 2548
rect 131236 2492 131246 2548
rect 134082 2492 134092 2548
rect 134148 2492 148316 2548
rect 148372 2492 148382 2548
rect 36754 2380 36764 2436
rect 36820 2380 83804 2436
rect 83860 2380 83870 2436
rect 91858 2380 91868 2436
rect 91924 2380 135996 2436
rect 136052 2380 136062 2436
rect 139682 2380 139692 2436
rect 139748 2380 166460 2436
rect 166516 2380 166526 2436
rect 110786 2268 110796 2324
rect 110852 2268 127820 2324
rect 127876 2268 127886 2324
rect 130722 2268 130732 2324
rect 130788 2268 162540 2324
rect 162596 2268 162606 2324
rect 105074 2156 105084 2212
rect 105140 2156 114716 2212
rect 114772 2156 114782 2212
rect 21634 1596 21644 1652
rect 21700 1596 79884 1652
rect 79940 1596 79950 1652
rect 97682 1596 97692 1652
rect 97748 1596 98588 1652
rect 98644 1596 98654 1652
rect 136098 1596 136108 1652
rect 136164 1596 169036 1652
rect 169092 1596 169102 1652
rect 60722 1484 60732 1540
rect 60788 1484 84812 1540
rect 84868 1484 84878 1540
rect 126802 1484 126812 1540
rect 126868 1484 155596 1540
rect 155652 1484 155662 1540
rect 35858 1372 35868 1428
rect 35924 1372 89292 1428
rect 89348 1372 89358 1428
rect 100482 1372 100492 1428
rect 100548 1372 111804 1428
rect 111860 1372 111870 1428
rect 114482 1372 114492 1428
rect 114548 1372 158620 1428
rect 158676 1372 158686 1428
rect 30818 1260 30828 1316
rect 30884 1260 82012 1316
rect 82068 1260 82078 1316
rect 123218 1260 123228 1316
rect 123284 1260 147756 1316
rect 147812 1260 147822 1316
rect 21746 1148 21756 1204
rect 21812 1148 70700 1204
rect 70756 1148 70766 1204
rect 126242 1148 126252 1204
rect 126308 1148 153468 1204
rect 153524 1148 153534 1204
rect 24770 1036 24780 1092
rect 24836 1036 64652 1092
rect 64708 1036 64718 1092
rect 85698 1036 85708 1092
rect 85764 1036 90748 1092
rect 129378 1036 129388 1092
rect 129444 1036 143388 1092
rect 143444 1036 143454 1092
rect 90692 980 90748 1036
rect 8306 924 8316 980
rect 8372 924 64092 980
rect 64148 924 64158 980
rect 87602 924 87612 980
rect 87668 924 87678 980
rect 90692 924 137676 980
rect 137732 924 137742 980
rect 87612 868 87668 924
rect 87612 812 140700 868
rect 140756 812 140766 868
rect 98578 700 98588 756
rect 98644 700 130508 756
rect 130564 700 130574 756
<< via3 >>
rect 4476 116788 4532 116844
rect 4580 116788 4636 116844
rect 4684 116788 4740 116844
rect 35196 116788 35252 116844
rect 35300 116788 35356 116844
rect 35404 116788 35460 116844
rect 65916 116788 65972 116844
rect 66020 116788 66076 116844
rect 66124 116788 66180 116844
rect 96636 116788 96692 116844
rect 96740 116788 96796 116844
rect 96844 116788 96900 116844
rect 127356 116788 127412 116844
rect 127460 116788 127516 116844
rect 127564 116788 127620 116844
rect 158076 116788 158132 116844
rect 158180 116788 158236 116844
rect 158284 116788 158340 116844
rect 95340 116172 95396 116228
rect 19836 116004 19892 116060
rect 19940 116004 19996 116060
rect 20044 116004 20100 116060
rect 50556 116004 50612 116060
rect 50660 116004 50716 116060
rect 50764 116004 50820 116060
rect 81276 116004 81332 116060
rect 81380 116004 81436 116060
rect 81484 116004 81540 116060
rect 111996 116004 112052 116060
rect 112100 116004 112156 116060
rect 112204 116004 112260 116060
rect 142716 116004 142772 116060
rect 142820 116004 142876 116060
rect 142924 116004 142980 116060
rect 173436 116004 173492 116060
rect 173540 116004 173596 116060
rect 173644 116004 173700 116060
rect 4476 115220 4532 115276
rect 4580 115220 4636 115276
rect 4684 115220 4740 115276
rect 35196 115220 35252 115276
rect 35300 115220 35356 115276
rect 35404 115220 35460 115276
rect 65916 115220 65972 115276
rect 66020 115220 66076 115276
rect 66124 115220 66180 115276
rect 96636 115220 96692 115276
rect 96740 115220 96796 115276
rect 96844 115220 96900 115276
rect 127356 115220 127412 115276
rect 127460 115220 127516 115276
rect 127564 115220 127620 115276
rect 158076 115220 158132 115276
rect 158180 115220 158236 115276
rect 158284 115220 158340 115276
rect 19836 114436 19892 114492
rect 19940 114436 19996 114492
rect 20044 114436 20100 114492
rect 50556 114436 50612 114492
rect 50660 114436 50716 114492
rect 50764 114436 50820 114492
rect 81276 114436 81332 114492
rect 81380 114436 81436 114492
rect 81484 114436 81540 114492
rect 111996 114436 112052 114492
rect 112100 114436 112156 114492
rect 112204 114436 112260 114492
rect 142716 114436 142772 114492
rect 142820 114436 142876 114492
rect 142924 114436 142980 114492
rect 173436 114436 173492 114492
rect 173540 114436 173596 114492
rect 173644 114436 173700 114492
rect 4476 113652 4532 113708
rect 4580 113652 4636 113708
rect 4684 113652 4740 113708
rect 35196 113652 35252 113708
rect 35300 113652 35356 113708
rect 35404 113652 35460 113708
rect 65916 113652 65972 113708
rect 66020 113652 66076 113708
rect 66124 113652 66180 113708
rect 96636 113652 96692 113708
rect 96740 113652 96796 113708
rect 96844 113652 96900 113708
rect 127356 113652 127412 113708
rect 127460 113652 127516 113708
rect 127564 113652 127620 113708
rect 158076 113652 158132 113708
rect 158180 113652 158236 113708
rect 158284 113652 158340 113708
rect 19836 112868 19892 112924
rect 19940 112868 19996 112924
rect 20044 112868 20100 112924
rect 50556 112868 50612 112924
rect 50660 112868 50716 112924
rect 50764 112868 50820 112924
rect 81276 112868 81332 112924
rect 81380 112868 81436 112924
rect 81484 112868 81540 112924
rect 111996 112868 112052 112924
rect 112100 112868 112156 112924
rect 112204 112868 112260 112924
rect 142716 112868 142772 112924
rect 142820 112868 142876 112924
rect 142924 112868 142980 112924
rect 173436 112868 173492 112924
rect 173540 112868 173596 112924
rect 173644 112868 173700 112924
rect 4476 112084 4532 112140
rect 4580 112084 4636 112140
rect 4684 112084 4740 112140
rect 35196 112084 35252 112140
rect 35300 112084 35356 112140
rect 35404 112084 35460 112140
rect 65916 112084 65972 112140
rect 66020 112084 66076 112140
rect 66124 112084 66180 112140
rect 96636 112084 96692 112140
rect 96740 112084 96796 112140
rect 96844 112084 96900 112140
rect 127356 112084 127412 112140
rect 127460 112084 127516 112140
rect 127564 112084 127620 112140
rect 158076 112084 158132 112140
rect 158180 112084 158236 112140
rect 158284 112084 158340 112140
rect 19836 111300 19892 111356
rect 19940 111300 19996 111356
rect 20044 111300 20100 111356
rect 50556 111300 50612 111356
rect 50660 111300 50716 111356
rect 50764 111300 50820 111356
rect 81276 111300 81332 111356
rect 81380 111300 81436 111356
rect 81484 111300 81540 111356
rect 111996 111300 112052 111356
rect 112100 111300 112156 111356
rect 112204 111300 112260 111356
rect 142716 111300 142772 111356
rect 142820 111300 142876 111356
rect 142924 111300 142980 111356
rect 173436 111300 173492 111356
rect 173540 111300 173596 111356
rect 173644 111300 173700 111356
rect 4476 110516 4532 110572
rect 4580 110516 4636 110572
rect 4684 110516 4740 110572
rect 35196 110516 35252 110572
rect 35300 110516 35356 110572
rect 35404 110516 35460 110572
rect 65916 110516 65972 110572
rect 66020 110516 66076 110572
rect 66124 110516 66180 110572
rect 96636 110516 96692 110572
rect 96740 110516 96796 110572
rect 96844 110516 96900 110572
rect 127356 110516 127412 110572
rect 127460 110516 127516 110572
rect 127564 110516 127620 110572
rect 158076 110516 158132 110572
rect 158180 110516 158236 110572
rect 158284 110516 158340 110572
rect 19836 109732 19892 109788
rect 19940 109732 19996 109788
rect 20044 109732 20100 109788
rect 50556 109732 50612 109788
rect 50660 109732 50716 109788
rect 50764 109732 50820 109788
rect 81276 109732 81332 109788
rect 81380 109732 81436 109788
rect 81484 109732 81540 109788
rect 111996 109732 112052 109788
rect 112100 109732 112156 109788
rect 112204 109732 112260 109788
rect 142716 109732 142772 109788
rect 142820 109732 142876 109788
rect 142924 109732 142980 109788
rect 173436 109732 173492 109788
rect 173540 109732 173596 109788
rect 173644 109732 173700 109788
rect 4476 108948 4532 109004
rect 4580 108948 4636 109004
rect 4684 108948 4740 109004
rect 35196 108948 35252 109004
rect 35300 108948 35356 109004
rect 35404 108948 35460 109004
rect 65916 108948 65972 109004
rect 66020 108948 66076 109004
rect 66124 108948 66180 109004
rect 96636 108948 96692 109004
rect 96740 108948 96796 109004
rect 96844 108948 96900 109004
rect 127356 108948 127412 109004
rect 127460 108948 127516 109004
rect 127564 108948 127620 109004
rect 158076 108948 158132 109004
rect 158180 108948 158236 109004
rect 158284 108948 158340 109004
rect 57148 108332 57204 108388
rect 19836 108164 19892 108220
rect 19940 108164 19996 108220
rect 20044 108164 20100 108220
rect 50556 108164 50612 108220
rect 50660 108164 50716 108220
rect 50764 108164 50820 108220
rect 81276 108164 81332 108220
rect 81380 108164 81436 108220
rect 81484 108164 81540 108220
rect 111996 108164 112052 108220
rect 112100 108164 112156 108220
rect 112204 108164 112260 108220
rect 142716 108164 142772 108220
rect 142820 108164 142876 108220
rect 142924 108164 142980 108220
rect 173436 108164 173492 108220
rect 173540 108164 173596 108220
rect 173644 108164 173700 108220
rect 4476 107380 4532 107436
rect 4580 107380 4636 107436
rect 4684 107380 4740 107436
rect 35196 107380 35252 107436
rect 35300 107380 35356 107436
rect 35404 107380 35460 107436
rect 65916 107380 65972 107436
rect 66020 107380 66076 107436
rect 66124 107380 66180 107436
rect 96636 107380 96692 107436
rect 96740 107380 96796 107436
rect 96844 107380 96900 107436
rect 127356 107380 127412 107436
rect 127460 107380 127516 107436
rect 127564 107380 127620 107436
rect 158076 107380 158132 107436
rect 158180 107380 158236 107436
rect 158284 107380 158340 107436
rect 19836 106596 19892 106652
rect 19940 106596 19996 106652
rect 20044 106596 20100 106652
rect 50556 106596 50612 106652
rect 50660 106596 50716 106652
rect 50764 106596 50820 106652
rect 81276 106596 81332 106652
rect 81380 106596 81436 106652
rect 81484 106596 81540 106652
rect 111996 106596 112052 106652
rect 112100 106596 112156 106652
rect 112204 106596 112260 106652
rect 142716 106596 142772 106652
rect 142820 106596 142876 106652
rect 142924 106596 142980 106652
rect 173436 106596 173492 106652
rect 173540 106596 173596 106652
rect 173644 106596 173700 106652
rect 4476 105812 4532 105868
rect 4580 105812 4636 105868
rect 4684 105812 4740 105868
rect 35196 105812 35252 105868
rect 35300 105812 35356 105868
rect 35404 105812 35460 105868
rect 65916 105812 65972 105868
rect 66020 105812 66076 105868
rect 66124 105812 66180 105868
rect 96636 105812 96692 105868
rect 96740 105812 96796 105868
rect 96844 105812 96900 105868
rect 127356 105812 127412 105868
rect 127460 105812 127516 105868
rect 127564 105812 127620 105868
rect 158076 105812 158132 105868
rect 158180 105812 158236 105868
rect 158284 105812 158340 105868
rect 19836 105028 19892 105084
rect 19940 105028 19996 105084
rect 20044 105028 20100 105084
rect 50556 105028 50612 105084
rect 50660 105028 50716 105084
rect 50764 105028 50820 105084
rect 81276 105028 81332 105084
rect 81380 105028 81436 105084
rect 81484 105028 81540 105084
rect 111996 105028 112052 105084
rect 112100 105028 112156 105084
rect 112204 105028 112260 105084
rect 142716 105028 142772 105084
rect 142820 105028 142876 105084
rect 142924 105028 142980 105084
rect 173436 105028 173492 105084
rect 173540 105028 173596 105084
rect 173644 105028 173700 105084
rect 4476 104244 4532 104300
rect 4580 104244 4636 104300
rect 4684 104244 4740 104300
rect 35196 104244 35252 104300
rect 35300 104244 35356 104300
rect 35404 104244 35460 104300
rect 65916 104244 65972 104300
rect 66020 104244 66076 104300
rect 66124 104244 66180 104300
rect 96636 104244 96692 104300
rect 96740 104244 96796 104300
rect 96844 104244 96900 104300
rect 127356 104244 127412 104300
rect 127460 104244 127516 104300
rect 127564 104244 127620 104300
rect 158076 104244 158132 104300
rect 158180 104244 158236 104300
rect 158284 104244 158340 104300
rect 19836 103460 19892 103516
rect 19940 103460 19996 103516
rect 20044 103460 20100 103516
rect 50556 103460 50612 103516
rect 50660 103460 50716 103516
rect 50764 103460 50820 103516
rect 81276 103460 81332 103516
rect 81380 103460 81436 103516
rect 81484 103460 81540 103516
rect 111996 103460 112052 103516
rect 112100 103460 112156 103516
rect 112204 103460 112260 103516
rect 142716 103460 142772 103516
rect 142820 103460 142876 103516
rect 142924 103460 142980 103516
rect 173436 103460 173492 103516
rect 173540 103460 173596 103516
rect 173644 103460 173700 103516
rect 4476 102676 4532 102732
rect 4580 102676 4636 102732
rect 4684 102676 4740 102732
rect 35196 102676 35252 102732
rect 35300 102676 35356 102732
rect 35404 102676 35460 102732
rect 65916 102676 65972 102732
rect 66020 102676 66076 102732
rect 66124 102676 66180 102732
rect 96636 102676 96692 102732
rect 96740 102676 96796 102732
rect 96844 102676 96900 102732
rect 127356 102676 127412 102732
rect 127460 102676 127516 102732
rect 127564 102676 127620 102732
rect 158076 102676 158132 102732
rect 158180 102676 158236 102732
rect 158284 102676 158340 102732
rect 19836 101892 19892 101948
rect 19940 101892 19996 101948
rect 20044 101892 20100 101948
rect 50556 101892 50612 101948
rect 50660 101892 50716 101948
rect 50764 101892 50820 101948
rect 81276 101892 81332 101948
rect 81380 101892 81436 101948
rect 81484 101892 81540 101948
rect 111996 101892 112052 101948
rect 112100 101892 112156 101948
rect 112204 101892 112260 101948
rect 142716 101892 142772 101948
rect 142820 101892 142876 101948
rect 142924 101892 142980 101948
rect 173436 101892 173492 101948
rect 173540 101892 173596 101948
rect 173644 101892 173700 101948
rect 4476 101108 4532 101164
rect 4580 101108 4636 101164
rect 4684 101108 4740 101164
rect 35196 101108 35252 101164
rect 35300 101108 35356 101164
rect 35404 101108 35460 101164
rect 65916 101108 65972 101164
rect 66020 101108 66076 101164
rect 66124 101108 66180 101164
rect 96636 101108 96692 101164
rect 96740 101108 96796 101164
rect 96844 101108 96900 101164
rect 127356 101108 127412 101164
rect 127460 101108 127516 101164
rect 127564 101108 127620 101164
rect 158076 101108 158132 101164
rect 158180 101108 158236 101164
rect 158284 101108 158340 101164
rect 19836 100324 19892 100380
rect 19940 100324 19996 100380
rect 20044 100324 20100 100380
rect 50556 100324 50612 100380
rect 50660 100324 50716 100380
rect 50764 100324 50820 100380
rect 81276 100324 81332 100380
rect 81380 100324 81436 100380
rect 81484 100324 81540 100380
rect 111996 100324 112052 100380
rect 112100 100324 112156 100380
rect 112204 100324 112260 100380
rect 142716 100324 142772 100380
rect 142820 100324 142876 100380
rect 142924 100324 142980 100380
rect 173436 100324 173492 100380
rect 173540 100324 173596 100380
rect 173644 100324 173700 100380
rect 4476 99540 4532 99596
rect 4580 99540 4636 99596
rect 4684 99540 4740 99596
rect 35196 99540 35252 99596
rect 35300 99540 35356 99596
rect 35404 99540 35460 99596
rect 65916 99540 65972 99596
rect 66020 99540 66076 99596
rect 66124 99540 66180 99596
rect 96636 99540 96692 99596
rect 96740 99540 96796 99596
rect 96844 99540 96900 99596
rect 127356 99540 127412 99596
rect 127460 99540 127516 99596
rect 127564 99540 127620 99596
rect 158076 99540 158132 99596
rect 158180 99540 158236 99596
rect 158284 99540 158340 99596
rect 19836 98756 19892 98812
rect 19940 98756 19996 98812
rect 20044 98756 20100 98812
rect 50556 98756 50612 98812
rect 50660 98756 50716 98812
rect 50764 98756 50820 98812
rect 81276 98756 81332 98812
rect 81380 98756 81436 98812
rect 81484 98756 81540 98812
rect 111996 98756 112052 98812
rect 112100 98756 112156 98812
rect 112204 98756 112260 98812
rect 142716 98756 142772 98812
rect 142820 98756 142876 98812
rect 142924 98756 142980 98812
rect 173436 98756 173492 98812
rect 173540 98756 173596 98812
rect 173644 98756 173700 98812
rect 4476 97972 4532 98028
rect 4580 97972 4636 98028
rect 4684 97972 4740 98028
rect 35196 97972 35252 98028
rect 35300 97972 35356 98028
rect 35404 97972 35460 98028
rect 65916 97972 65972 98028
rect 66020 97972 66076 98028
rect 66124 97972 66180 98028
rect 96636 97972 96692 98028
rect 96740 97972 96796 98028
rect 96844 97972 96900 98028
rect 127356 97972 127412 98028
rect 127460 97972 127516 98028
rect 127564 97972 127620 98028
rect 158076 97972 158132 98028
rect 158180 97972 158236 98028
rect 158284 97972 158340 98028
rect 19836 97188 19892 97244
rect 19940 97188 19996 97244
rect 20044 97188 20100 97244
rect 50556 97188 50612 97244
rect 50660 97188 50716 97244
rect 50764 97188 50820 97244
rect 81276 97188 81332 97244
rect 81380 97188 81436 97244
rect 81484 97188 81540 97244
rect 111996 97188 112052 97244
rect 112100 97188 112156 97244
rect 112204 97188 112260 97244
rect 142716 97188 142772 97244
rect 142820 97188 142876 97244
rect 142924 97188 142980 97244
rect 173436 97188 173492 97244
rect 173540 97188 173596 97244
rect 173644 97188 173700 97244
rect 4476 96404 4532 96460
rect 4580 96404 4636 96460
rect 4684 96404 4740 96460
rect 35196 96404 35252 96460
rect 35300 96404 35356 96460
rect 35404 96404 35460 96460
rect 65916 96404 65972 96460
rect 66020 96404 66076 96460
rect 66124 96404 66180 96460
rect 96636 96404 96692 96460
rect 96740 96404 96796 96460
rect 96844 96404 96900 96460
rect 127356 96404 127412 96460
rect 127460 96404 127516 96460
rect 127564 96404 127620 96460
rect 158076 96404 158132 96460
rect 158180 96404 158236 96460
rect 158284 96404 158340 96460
rect 19836 95620 19892 95676
rect 19940 95620 19996 95676
rect 20044 95620 20100 95676
rect 50556 95620 50612 95676
rect 50660 95620 50716 95676
rect 50764 95620 50820 95676
rect 81276 95620 81332 95676
rect 81380 95620 81436 95676
rect 81484 95620 81540 95676
rect 111996 95620 112052 95676
rect 112100 95620 112156 95676
rect 112204 95620 112260 95676
rect 142716 95620 142772 95676
rect 142820 95620 142876 95676
rect 142924 95620 142980 95676
rect 173436 95620 173492 95676
rect 173540 95620 173596 95676
rect 173644 95620 173700 95676
rect 4476 94836 4532 94892
rect 4580 94836 4636 94892
rect 4684 94836 4740 94892
rect 35196 94836 35252 94892
rect 35300 94836 35356 94892
rect 35404 94836 35460 94892
rect 65916 94836 65972 94892
rect 66020 94836 66076 94892
rect 66124 94836 66180 94892
rect 96636 94836 96692 94892
rect 96740 94836 96796 94892
rect 96844 94836 96900 94892
rect 127356 94836 127412 94892
rect 127460 94836 127516 94892
rect 127564 94836 127620 94892
rect 158076 94836 158132 94892
rect 158180 94836 158236 94892
rect 158284 94836 158340 94892
rect 19836 94052 19892 94108
rect 19940 94052 19996 94108
rect 20044 94052 20100 94108
rect 50556 94052 50612 94108
rect 50660 94052 50716 94108
rect 50764 94052 50820 94108
rect 81276 94052 81332 94108
rect 81380 94052 81436 94108
rect 81484 94052 81540 94108
rect 111996 94052 112052 94108
rect 112100 94052 112156 94108
rect 112204 94052 112260 94108
rect 142716 94052 142772 94108
rect 142820 94052 142876 94108
rect 142924 94052 142980 94108
rect 173436 94052 173492 94108
rect 173540 94052 173596 94108
rect 173644 94052 173700 94108
rect 4476 93268 4532 93324
rect 4580 93268 4636 93324
rect 4684 93268 4740 93324
rect 35196 93268 35252 93324
rect 35300 93268 35356 93324
rect 35404 93268 35460 93324
rect 65916 93268 65972 93324
rect 66020 93268 66076 93324
rect 66124 93268 66180 93324
rect 96636 93268 96692 93324
rect 96740 93268 96796 93324
rect 96844 93268 96900 93324
rect 127356 93268 127412 93324
rect 127460 93268 127516 93324
rect 127564 93268 127620 93324
rect 158076 93268 158132 93324
rect 158180 93268 158236 93324
rect 158284 93268 158340 93324
rect 19836 92484 19892 92540
rect 19940 92484 19996 92540
rect 20044 92484 20100 92540
rect 50556 92484 50612 92540
rect 50660 92484 50716 92540
rect 50764 92484 50820 92540
rect 81276 92484 81332 92540
rect 81380 92484 81436 92540
rect 81484 92484 81540 92540
rect 111996 92484 112052 92540
rect 112100 92484 112156 92540
rect 112204 92484 112260 92540
rect 142716 92484 142772 92540
rect 142820 92484 142876 92540
rect 142924 92484 142980 92540
rect 173436 92484 173492 92540
rect 173540 92484 173596 92540
rect 173644 92484 173700 92540
rect 4476 91700 4532 91756
rect 4580 91700 4636 91756
rect 4684 91700 4740 91756
rect 35196 91700 35252 91756
rect 35300 91700 35356 91756
rect 35404 91700 35460 91756
rect 65916 91700 65972 91756
rect 66020 91700 66076 91756
rect 66124 91700 66180 91756
rect 96636 91700 96692 91756
rect 96740 91700 96796 91756
rect 96844 91700 96900 91756
rect 127356 91700 127412 91756
rect 127460 91700 127516 91756
rect 127564 91700 127620 91756
rect 158076 91700 158132 91756
rect 158180 91700 158236 91756
rect 158284 91700 158340 91756
rect 19836 90916 19892 90972
rect 19940 90916 19996 90972
rect 20044 90916 20100 90972
rect 50556 90916 50612 90972
rect 50660 90916 50716 90972
rect 50764 90916 50820 90972
rect 81276 90916 81332 90972
rect 81380 90916 81436 90972
rect 81484 90916 81540 90972
rect 111996 90916 112052 90972
rect 112100 90916 112156 90972
rect 112204 90916 112260 90972
rect 142716 90916 142772 90972
rect 142820 90916 142876 90972
rect 142924 90916 142980 90972
rect 173436 90916 173492 90972
rect 173540 90916 173596 90972
rect 173644 90916 173700 90972
rect 4476 90132 4532 90188
rect 4580 90132 4636 90188
rect 4684 90132 4740 90188
rect 35196 90132 35252 90188
rect 35300 90132 35356 90188
rect 35404 90132 35460 90188
rect 65916 90132 65972 90188
rect 66020 90132 66076 90188
rect 66124 90132 66180 90188
rect 96636 90132 96692 90188
rect 96740 90132 96796 90188
rect 96844 90132 96900 90188
rect 127356 90132 127412 90188
rect 127460 90132 127516 90188
rect 127564 90132 127620 90188
rect 158076 90132 158132 90188
rect 158180 90132 158236 90188
rect 158284 90132 158340 90188
rect 19836 89348 19892 89404
rect 19940 89348 19996 89404
rect 20044 89348 20100 89404
rect 50556 89348 50612 89404
rect 50660 89348 50716 89404
rect 50764 89348 50820 89404
rect 81276 89348 81332 89404
rect 81380 89348 81436 89404
rect 81484 89348 81540 89404
rect 111996 89348 112052 89404
rect 112100 89348 112156 89404
rect 112204 89348 112260 89404
rect 142716 89348 142772 89404
rect 142820 89348 142876 89404
rect 142924 89348 142980 89404
rect 173436 89348 173492 89404
rect 173540 89348 173596 89404
rect 173644 89348 173700 89404
rect 4476 88564 4532 88620
rect 4580 88564 4636 88620
rect 4684 88564 4740 88620
rect 35196 88564 35252 88620
rect 35300 88564 35356 88620
rect 35404 88564 35460 88620
rect 65916 88564 65972 88620
rect 66020 88564 66076 88620
rect 66124 88564 66180 88620
rect 96636 88564 96692 88620
rect 96740 88564 96796 88620
rect 96844 88564 96900 88620
rect 127356 88564 127412 88620
rect 127460 88564 127516 88620
rect 127564 88564 127620 88620
rect 158076 88564 158132 88620
rect 158180 88564 158236 88620
rect 158284 88564 158340 88620
rect 19836 87780 19892 87836
rect 19940 87780 19996 87836
rect 20044 87780 20100 87836
rect 50556 87780 50612 87836
rect 50660 87780 50716 87836
rect 50764 87780 50820 87836
rect 81276 87780 81332 87836
rect 81380 87780 81436 87836
rect 81484 87780 81540 87836
rect 111996 87780 112052 87836
rect 112100 87780 112156 87836
rect 112204 87780 112260 87836
rect 142716 87780 142772 87836
rect 142820 87780 142876 87836
rect 142924 87780 142980 87836
rect 173436 87780 173492 87836
rect 173540 87780 173596 87836
rect 173644 87780 173700 87836
rect 4476 86996 4532 87052
rect 4580 86996 4636 87052
rect 4684 86996 4740 87052
rect 35196 86996 35252 87052
rect 35300 86996 35356 87052
rect 35404 86996 35460 87052
rect 65916 86996 65972 87052
rect 66020 86996 66076 87052
rect 66124 86996 66180 87052
rect 96636 86996 96692 87052
rect 96740 86996 96796 87052
rect 96844 86996 96900 87052
rect 127356 86996 127412 87052
rect 127460 86996 127516 87052
rect 127564 86996 127620 87052
rect 158076 86996 158132 87052
rect 158180 86996 158236 87052
rect 158284 86996 158340 87052
rect 19836 86212 19892 86268
rect 19940 86212 19996 86268
rect 20044 86212 20100 86268
rect 50556 86212 50612 86268
rect 50660 86212 50716 86268
rect 50764 86212 50820 86268
rect 81276 86212 81332 86268
rect 81380 86212 81436 86268
rect 81484 86212 81540 86268
rect 111996 86212 112052 86268
rect 112100 86212 112156 86268
rect 112204 86212 112260 86268
rect 142716 86212 142772 86268
rect 142820 86212 142876 86268
rect 142924 86212 142980 86268
rect 173436 86212 173492 86268
rect 173540 86212 173596 86268
rect 173644 86212 173700 86268
rect 4476 85428 4532 85484
rect 4580 85428 4636 85484
rect 4684 85428 4740 85484
rect 35196 85428 35252 85484
rect 35300 85428 35356 85484
rect 35404 85428 35460 85484
rect 65916 85428 65972 85484
rect 66020 85428 66076 85484
rect 66124 85428 66180 85484
rect 96636 85428 96692 85484
rect 96740 85428 96796 85484
rect 96844 85428 96900 85484
rect 127356 85428 127412 85484
rect 127460 85428 127516 85484
rect 127564 85428 127620 85484
rect 158076 85428 158132 85484
rect 158180 85428 158236 85484
rect 158284 85428 158340 85484
rect 19836 84644 19892 84700
rect 19940 84644 19996 84700
rect 20044 84644 20100 84700
rect 50556 84644 50612 84700
rect 50660 84644 50716 84700
rect 50764 84644 50820 84700
rect 81276 84644 81332 84700
rect 81380 84644 81436 84700
rect 81484 84644 81540 84700
rect 111996 84644 112052 84700
rect 112100 84644 112156 84700
rect 112204 84644 112260 84700
rect 142716 84644 142772 84700
rect 142820 84644 142876 84700
rect 142924 84644 142980 84700
rect 173436 84644 173492 84700
rect 173540 84644 173596 84700
rect 173644 84644 173700 84700
rect 4476 83860 4532 83916
rect 4580 83860 4636 83916
rect 4684 83860 4740 83916
rect 35196 83860 35252 83916
rect 35300 83860 35356 83916
rect 35404 83860 35460 83916
rect 65916 83860 65972 83916
rect 66020 83860 66076 83916
rect 66124 83860 66180 83916
rect 96636 83860 96692 83916
rect 96740 83860 96796 83916
rect 96844 83860 96900 83916
rect 127356 83860 127412 83916
rect 127460 83860 127516 83916
rect 127564 83860 127620 83916
rect 158076 83860 158132 83916
rect 158180 83860 158236 83916
rect 158284 83860 158340 83916
rect 19836 83076 19892 83132
rect 19940 83076 19996 83132
rect 20044 83076 20100 83132
rect 50556 83076 50612 83132
rect 50660 83076 50716 83132
rect 50764 83076 50820 83132
rect 81276 83076 81332 83132
rect 81380 83076 81436 83132
rect 81484 83076 81540 83132
rect 111996 83076 112052 83132
rect 112100 83076 112156 83132
rect 112204 83076 112260 83132
rect 142716 83076 142772 83132
rect 142820 83076 142876 83132
rect 142924 83076 142980 83132
rect 173436 83076 173492 83132
rect 173540 83076 173596 83132
rect 173644 83076 173700 83132
rect 4476 82292 4532 82348
rect 4580 82292 4636 82348
rect 4684 82292 4740 82348
rect 35196 82292 35252 82348
rect 35300 82292 35356 82348
rect 35404 82292 35460 82348
rect 65916 82292 65972 82348
rect 66020 82292 66076 82348
rect 66124 82292 66180 82348
rect 96636 82292 96692 82348
rect 96740 82292 96796 82348
rect 96844 82292 96900 82348
rect 127356 82292 127412 82348
rect 127460 82292 127516 82348
rect 127564 82292 127620 82348
rect 158076 82292 158132 82348
rect 158180 82292 158236 82348
rect 158284 82292 158340 82348
rect 19836 81508 19892 81564
rect 19940 81508 19996 81564
rect 20044 81508 20100 81564
rect 50556 81508 50612 81564
rect 50660 81508 50716 81564
rect 50764 81508 50820 81564
rect 81276 81508 81332 81564
rect 81380 81508 81436 81564
rect 81484 81508 81540 81564
rect 111996 81508 112052 81564
rect 112100 81508 112156 81564
rect 112204 81508 112260 81564
rect 142716 81508 142772 81564
rect 142820 81508 142876 81564
rect 142924 81508 142980 81564
rect 173436 81508 173492 81564
rect 173540 81508 173596 81564
rect 173644 81508 173700 81564
rect 4476 80724 4532 80780
rect 4580 80724 4636 80780
rect 4684 80724 4740 80780
rect 35196 80724 35252 80780
rect 35300 80724 35356 80780
rect 35404 80724 35460 80780
rect 65916 80724 65972 80780
rect 66020 80724 66076 80780
rect 66124 80724 66180 80780
rect 96636 80724 96692 80780
rect 96740 80724 96796 80780
rect 96844 80724 96900 80780
rect 127356 80724 127412 80780
rect 127460 80724 127516 80780
rect 127564 80724 127620 80780
rect 158076 80724 158132 80780
rect 158180 80724 158236 80780
rect 158284 80724 158340 80780
rect 19836 79940 19892 79996
rect 19940 79940 19996 79996
rect 20044 79940 20100 79996
rect 50556 79940 50612 79996
rect 50660 79940 50716 79996
rect 50764 79940 50820 79996
rect 81276 79940 81332 79996
rect 81380 79940 81436 79996
rect 81484 79940 81540 79996
rect 111996 79940 112052 79996
rect 112100 79940 112156 79996
rect 112204 79940 112260 79996
rect 142716 79940 142772 79996
rect 142820 79940 142876 79996
rect 142924 79940 142980 79996
rect 173436 79940 173492 79996
rect 173540 79940 173596 79996
rect 173644 79940 173700 79996
rect 4476 79156 4532 79212
rect 4580 79156 4636 79212
rect 4684 79156 4740 79212
rect 35196 79156 35252 79212
rect 35300 79156 35356 79212
rect 35404 79156 35460 79212
rect 65916 79156 65972 79212
rect 66020 79156 66076 79212
rect 66124 79156 66180 79212
rect 96636 79156 96692 79212
rect 96740 79156 96796 79212
rect 96844 79156 96900 79212
rect 127356 79156 127412 79212
rect 127460 79156 127516 79212
rect 127564 79156 127620 79212
rect 158076 79156 158132 79212
rect 158180 79156 158236 79212
rect 158284 79156 158340 79212
rect 19836 78372 19892 78428
rect 19940 78372 19996 78428
rect 20044 78372 20100 78428
rect 50556 78372 50612 78428
rect 50660 78372 50716 78428
rect 50764 78372 50820 78428
rect 81276 78372 81332 78428
rect 81380 78372 81436 78428
rect 81484 78372 81540 78428
rect 111996 78372 112052 78428
rect 112100 78372 112156 78428
rect 112204 78372 112260 78428
rect 142716 78372 142772 78428
rect 142820 78372 142876 78428
rect 142924 78372 142980 78428
rect 173436 78372 173492 78428
rect 173540 78372 173596 78428
rect 173644 78372 173700 78428
rect 4476 77588 4532 77644
rect 4580 77588 4636 77644
rect 4684 77588 4740 77644
rect 35196 77588 35252 77644
rect 35300 77588 35356 77644
rect 35404 77588 35460 77644
rect 65916 77588 65972 77644
rect 66020 77588 66076 77644
rect 66124 77588 66180 77644
rect 96636 77588 96692 77644
rect 96740 77588 96796 77644
rect 96844 77588 96900 77644
rect 127356 77588 127412 77644
rect 127460 77588 127516 77644
rect 127564 77588 127620 77644
rect 158076 77588 158132 77644
rect 158180 77588 158236 77644
rect 158284 77588 158340 77644
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 81276 76804 81332 76860
rect 81380 76804 81436 76860
rect 81484 76804 81540 76860
rect 111996 76804 112052 76860
rect 112100 76804 112156 76860
rect 112204 76804 112260 76860
rect 142716 76804 142772 76860
rect 142820 76804 142876 76860
rect 142924 76804 142980 76860
rect 173436 76804 173492 76860
rect 173540 76804 173596 76860
rect 173644 76804 173700 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 96636 76020 96692 76076
rect 96740 76020 96796 76076
rect 96844 76020 96900 76076
rect 127356 76020 127412 76076
rect 127460 76020 127516 76076
rect 127564 76020 127620 76076
rect 158076 76020 158132 76076
rect 158180 76020 158236 76076
rect 158284 76020 158340 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 81276 75236 81332 75292
rect 81380 75236 81436 75292
rect 81484 75236 81540 75292
rect 111996 75236 112052 75292
rect 112100 75236 112156 75292
rect 112204 75236 112260 75292
rect 142716 75236 142772 75292
rect 142820 75236 142876 75292
rect 142924 75236 142980 75292
rect 173436 75236 173492 75292
rect 173540 75236 173596 75292
rect 173644 75236 173700 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 96636 74452 96692 74508
rect 96740 74452 96796 74508
rect 96844 74452 96900 74508
rect 127356 74452 127412 74508
rect 127460 74452 127516 74508
rect 127564 74452 127620 74508
rect 158076 74452 158132 74508
rect 158180 74452 158236 74508
rect 158284 74452 158340 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 81276 73668 81332 73724
rect 81380 73668 81436 73724
rect 81484 73668 81540 73724
rect 111996 73668 112052 73724
rect 112100 73668 112156 73724
rect 112204 73668 112260 73724
rect 142716 73668 142772 73724
rect 142820 73668 142876 73724
rect 142924 73668 142980 73724
rect 173436 73668 173492 73724
rect 173540 73668 173596 73724
rect 173644 73668 173700 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 96636 72884 96692 72940
rect 96740 72884 96796 72940
rect 96844 72884 96900 72940
rect 127356 72884 127412 72940
rect 127460 72884 127516 72940
rect 127564 72884 127620 72940
rect 158076 72884 158132 72940
rect 158180 72884 158236 72940
rect 158284 72884 158340 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 81276 72100 81332 72156
rect 81380 72100 81436 72156
rect 81484 72100 81540 72156
rect 111996 72100 112052 72156
rect 112100 72100 112156 72156
rect 112204 72100 112260 72156
rect 142716 72100 142772 72156
rect 142820 72100 142876 72156
rect 142924 72100 142980 72156
rect 173436 72100 173492 72156
rect 173540 72100 173596 72156
rect 173644 72100 173700 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 96636 71316 96692 71372
rect 96740 71316 96796 71372
rect 96844 71316 96900 71372
rect 127356 71316 127412 71372
rect 127460 71316 127516 71372
rect 127564 71316 127620 71372
rect 158076 71316 158132 71372
rect 158180 71316 158236 71372
rect 158284 71316 158340 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 81276 70532 81332 70588
rect 81380 70532 81436 70588
rect 81484 70532 81540 70588
rect 111996 70532 112052 70588
rect 112100 70532 112156 70588
rect 112204 70532 112260 70588
rect 142716 70532 142772 70588
rect 142820 70532 142876 70588
rect 142924 70532 142980 70588
rect 173436 70532 173492 70588
rect 173540 70532 173596 70588
rect 173644 70532 173700 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 96636 69748 96692 69804
rect 96740 69748 96796 69804
rect 96844 69748 96900 69804
rect 127356 69748 127412 69804
rect 127460 69748 127516 69804
rect 127564 69748 127620 69804
rect 158076 69748 158132 69804
rect 158180 69748 158236 69804
rect 158284 69748 158340 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 81276 68964 81332 69020
rect 81380 68964 81436 69020
rect 81484 68964 81540 69020
rect 111996 68964 112052 69020
rect 112100 68964 112156 69020
rect 112204 68964 112260 69020
rect 142716 68964 142772 69020
rect 142820 68964 142876 69020
rect 142924 68964 142980 69020
rect 173436 68964 173492 69020
rect 173540 68964 173596 69020
rect 173644 68964 173700 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 96636 68180 96692 68236
rect 96740 68180 96796 68236
rect 96844 68180 96900 68236
rect 127356 68180 127412 68236
rect 127460 68180 127516 68236
rect 127564 68180 127620 68236
rect 158076 68180 158132 68236
rect 158180 68180 158236 68236
rect 158284 68180 158340 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 81276 67396 81332 67452
rect 81380 67396 81436 67452
rect 81484 67396 81540 67452
rect 111996 67396 112052 67452
rect 112100 67396 112156 67452
rect 112204 67396 112260 67452
rect 142716 67396 142772 67452
rect 142820 67396 142876 67452
rect 142924 67396 142980 67452
rect 173436 67396 173492 67452
rect 173540 67396 173596 67452
rect 173644 67396 173700 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 96636 66612 96692 66668
rect 96740 66612 96796 66668
rect 96844 66612 96900 66668
rect 127356 66612 127412 66668
rect 127460 66612 127516 66668
rect 127564 66612 127620 66668
rect 158076 66612 158132 66668
rect 158180 66612 158236 66668
rect 158284 66612 158340 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 81276 65828 81332 65884
rect 81380 65828 81436 65884
rect 81484 65828 81540 65884
rect 111996 65828 112052 65884
rect 112100 65828 112156 65884
rect 112204 65828 112260 65884
rect 142716 65828 142772 65884
rect 142820 65828 142876 65884
rect 142924 65828 142980 65884
rect 173436 65828 173492 65884
rect 173540 65828 173596 65884
rect 173644 65828 173700 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 96636 65044 96692 65100
rect 96740 65044 96796 65100
rect 96844 65044 96900 65100
rect 127356 65044 127412 65100
rect 127460 65044 127516 65100
rect 127564 65044 127620 65100
rect 158076 65044 158132 65100
rect 158180 65044 158236 65100
rect 158284 65044 158340 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 81276 64260 81332 64316
rect 81380 64260 81436 64316
rect 81484 64260 81540 64316
rect 111996 64260 112052 64316
rect 112100 64260 112156 64316
rect 112204 64260 112260 64316
rect 142716 64260 142772 64316
rect 142820 64260 142876 64316
rect 142924 64260 142980 64316
rect 173436 64260 173492 64316
rect 173540 64260 173596 64316
rect 173644 64260 173700 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 96636 63476 96692 63532
rect 96740 63476 96796 63532
rect 96844 63476 96900 63532
rect 127356 63476 127412 63532
rect 127460 63476 127516 63532
rect 127564 63476 127620 63532
rect 158076 63476 158132 63532
rect 158180 63476 158236 63532
rect 158284 63476 158340 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 81276 62692 81332 62748
rect 81380 62692 81436 62748
rect 81484 62692 81540 62748
rect 111996 62692 112052 62748
rect 112100 62692 112156 62748
rect 112204 62692 112260 62748
rect 142716 62692 142772 62748
rect 142820 62692 142876 62748
rect 142924 62692 142980 62748
rect 173436 62692 173492 62748
rect 173540 62692 173596 62748
rect 173644 62692 173700 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 96636 61908 96692 61964
rect 96740 61908 96796 61964
rect 96844 61908 96900 61964
rect 127356 61908 127412 61964
rect 127460 61908 127516 61964
rect 127564 61908 127620 61964
rect 158076 61908 158132 61964
rect 158180 61908 158236 61964
rect 158284 61908 158340 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 81276 61124 81332 61180
rect 81380 61124 81436 61180
rect 81484 61124 81540 61180
rect 111996 61124 112052 61180
rect 112100 61124 112156 61180
rect 112204 61124 112260 61180
rect 142716 61124 142772 61180
rect 142820 61124 142876 61180
rect 142924 61124 142980 61180
rect 173436 61124 173492 61180
rect 173540 61124 173596 61180
rect 173644 61124 173700 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 96636 60340 96692 60396
rect 96740 60340 96796 60396
rect 96844 60340 96900 60396
rect 127356 60340 127412 60396
rect 127460 60340 127516 60396
rect 127564 60340 127620 60396
rect 158076 60340 158132 60396
rect 158180 60340 158236 60396
rect 158284 60340 158340 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 81276 59556 81332 59612
rect 81380 59556 81436 59612
rect 81484 59556 81540 59612
rect 111996 59556 112052 59612
rect 112100 59556 112156 59612
rect 112204 59556 112260 59612
rect 142716 59556 142772 59612
rect 142820 59556 142876 59612
rect 142924 59556 142980 59612
rect 173436 59556 173492 59612
rect 173540 59556 173596 59612
rect 173644 59556 173700 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 96636 58772 96692 58828
rect 96740 58772 96796 58828
rect 96844 58772 96900 58828
rect 127356 58772 127412 58828
rect 127460 58772 127516 58828
rect 127564 58772 127620 58828
rect 158076 58772 158132 58828
rect 158180 58772 158236 58828
rect 158284 58772 158340 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 81276 57988 81332 58044
rect 81380 57988 81436 58044
rect 81484 57988 81540 58044
rect 111996 57988 112052 58044
rect 112100 57988 112156 58044
rect 112204 57988 112260 58044
rect 142716 57988 142772 58044
rect 142820 57988 142876 58044
rect 142924 57988 142980 58044
rect 173436 57988 173492 58044
rect 173540 57988 173596 58044
rect 173644 57988 173700 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 96636 57204 96692 57260
rect 96740 57204 96796 57260
rect 96844 57204 96900 57260
rect 127356 57204 127412 57260
rect 127460 57204 127516 57260
rect 127564 57204 127620 57260
rect 158076 57204 158132 57260
rect 158180 57204 158236 57260
rect 158284 57204 158340 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 81276 56420 81332 56476
rect 81380 56420 81436 56476
rect 81484 56420 81540 56476
rect 111996 56420 112052 56476
rect 112100 56420 112156 56476
rect 112204 56420 112260 56476
rect 142716 56420 142772 56476
rect 142820 56420 142876 56476
rect 142924 56420 142980 56476
rect 173436 56420 173492 56476
rect 173540 56420 173596 56476
rect 173644 56420 173700 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 96636 55636 96692 55692
rect 96740 55636 96796 55692
rect 96844 55636 96900 55692
rect 127356 55636 127412 55692
rect 127460 55636 127516 55692
rect 127564 55636 127620 55692
rect 158076 55636 158132 55692
rect 158180 55636 158236 55692
rect 158284 55636 158340 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 81276 54852 81332 54908
rect 81380 54852 81436 54908
rect 81484 54852 81540 54908
rect 111996 54852 112052 54908
rect 112100 54852 112156 54908
rect 112204 54852 112260 54908
rect 142716 54852 142772 54908
rect 142820 54852 142876 54908
rect 142924 54852 142980 54908
rect 173436 54852 173492 54908
rect 173540 54852 173596 54908
rect 173644 54852 173700 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 96636 54068 96692 54124
rect 96740 54068 96796 54124
rect 96844 54068 96900 54124
rect 127356 54068 127412 54124
rect 127460 54068 127516 54124
rect 127564 54068 127620 54124
rect 158076 54068 158132 54124
rect 158180 54068 158236 54124
rect 158284 54068 158340 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 81276 53284 81332 53340
rect 81380 53284 81436 53340
rect 81484 53284 81540 53340
rect 111996 53284 112052 53340
rect 112100 53284 112156 53340
rect 112204 53284 112260 53340
rect 142716 53284 142772 53340
rect 142820 53284 142876 53340
rect 142924 53284 142980 53340
rect 173436 53284 173492 53340
rect 173540 53284 173596 53340
rect 173644 53284 173700 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 96636 52500 96692 52556
rect 96740 52500 96796 52556
rect 96844 52500 96900 52556
rect 127356 52500 127412 52556
rect 127460 52500 127516 52556
rect 127564 52500 127620 52556
rect 158076 52500 158132 52556
rect 158180 52500 158236 52556
rect 158284 52500 158340 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 81276 51716 81332 51772
rect 81380 51716 81436 51772
rect 81484 51716 81540 51772
rect 111996 51716 112052 51772
rect 112100 51716 112156 51772
rect 112204 51716 112260 51772
rect 142716 51716 142772 51772
rect 142820 51716 142876 51772
rect 142924 51716 142980 51772
rect 173436 51716 173492 51772
rect 173540 51716 173596 51772
rect 173644 51716 173700 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 96636 50932 96692 50988
rect 96740 50932 96796 50988
rect 96844 50932 96900 50988
rect 127356 50932 127412 50988
rect 127460 50932 127516 50988
rect 127564 50932 127620 50988
rect 158076 50932 158132 50988
rect 158180 50932 158236 50988
rect 158284 50932 158340 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 81276 50148 81332 50204
rect 81380 50148 81436 50204
rect 81484 50148 81540 50204
rect 111996 50148 112052 50204
rect 112100 50148 112156 50204
rect 112204 50148 112260 50204
rect 142716 50148 142772 50204
rect 142820 50148 142876 50204
rect 142924 50148 142980 50204
rect 173436 50148 173492 50204
rect 173540 50148 173596 50204
rect 173644 50148 173700 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 96636 49364 96692 49420
rect 96740 49364 96796 49420
rect 96844 49364 96900 49420
rect 127356 49364 127412 49420
rect 127460 49364 127516 49420
rect 127564 49364 127620 49420
rect 158076 49364 158132 49420
rect 158180 49364 158236 49420
rect 158284 49364 158340 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 81276 48580 81332 48636
rect 81380 48580 81436 48636
rect 81484 48580 81540 48636
rect 111996 48580 112052 48636
rect 112100 48580 112156 48636
rect 112204 48580 112260 48636
rect 142716 48580 142772 48636
rect 142820 48580 142876 48636
rect 142924 48580 142980 48636
rect 173436 48580 173492 48636
rect 173540 48580 173596 48636
rect 173644 48580 173700 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 96636 47796 96692 47852
rect 96740 47796 96796 47852
rect 96844 47796 96900 47852
rect 127356 47796 127412 47852
rect 127460 47796 127516 47852
rect 127564 47796 127620 47852
rect 158076 47796 158132 47852
rect 158180 47796 158236 47852
rect 158284 47796 158340 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 81276 47012 81332 47068
rect 81380 47012 81436 47068
rect 81484 47012 81540 47068
rect 111996 47012 112052 47068
rect 112100 47012 112156 47068
rect 112204 47012 112260 47068
rect 142716 47012 142772 47068
rect 142820 47012 142876 47068
rect 142924 47012 142980 47068
rect 173436 47012 173492 47068
rect 173540 47012 173596 47068
rect 173644 47012 173700 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 96636 46228 96692 46284
rect 96740 46228 96796 46284
rect 96844 46228 96900 46284
rect 127356 46228 127412 46284
rect 127460 46228 127516 46284
rect 127564 46228 127620 46284
rect 158076 46228 158132 46284
rect 158180 46228 158236 46284
rect 158284 46228 158340 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 81276 45444 81332 45500
rect 81380 45444 81436 45500
rect 81484 45444 81540 45500
rect 111996 45444 112052 45500
rect 112100 45444 112156 45500
rect 112204 45444 112260 45500
rect 142716 45444 142772 45500
rect 142820 45444 142876 45500
rect 142924 45444 142980 45500
rect 173436 45444 173492 45500
rect 173540 45444 173596 45500
rect 173644 45444 173700 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 96636 44660 96692 44716
rect 96740 44660 96796 44716
rect 96844 44660 96900 44716
rect 127356 44660 127412 44716
rect 127460 44660 127516 44716
rect 127564 44660 127620 44716
rect 158076 44660 158132 44716
rect 158180 44660 158236 44716
rect 158284 44660 158340 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 81276 43876 81332 43932
rect 81380 43876 81436 43932
rect 81484 43876 81540 43932
rect 111996 43876 112052 43932
rect 112100 43876 112156 43932
rect 112204 43876 112260 43932
rect 142716 43876 142772 43932
rect 142820 43876 142876 43932
rect 142924 43876 142980 43932
rect 173436 43876 173492 43932
rect 173540 43876 173596 43932
rect 173644 43876 173700 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 96636 43092 96692 43148
rect 96740 43092 96796 43148
rect 96844 43092 96900 43148
rect 127356 43092 127412 43148
rect 127460 43092 127516 43148
rect 127564 43092 127620 43148
rect 158076 43092 158132 43148
rect 158180 43092 158236 43148
rect 158284 43092 158340 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 81276 42308 81332 42364
rect 81380 42308 81436 42364
rect 81484 42308 81540 42364
rect 111996 42308 112052 42364
rect 112100 42308 112156 42364
rect 112204 42308 112260 42364
rect 142716 42308 142772 42364
rect 142820 42308 142876 42364
rect 142924 42308 142980 42364
rect 173436 42308 173492 42364
rect 173540 42308 173596 42364
rect 173644 42308 173700 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 96636 41524 96692 41580
rect 96740 41524 96796 41580
rect 96844 41524 96900 41580
rect 127356 41524 127412 41580
rect 127460 41524 127516 41580
rect 127564 41524 127620 41580
rect 158076 41524 158132 41580
rect 158180 41524 158236 41580
rect 158284 41524 158340 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 81276 40740 81332 40796
rect 81380 40740 81436 40796
rect 81484 40740 81540 40796
rect 111996 40740 112052 40796
rect 112100 40740 112156 40796
rect 112204 40740 112260 40796
rect 142716 40740 142772 40796
rect 142820 40740 142876 40796
rect 142924 40740 142980 40796
rect 173436 40740 173492 40796
rect 173540 40740 173596 40796
rect 173644 40740 173700 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 96636 39956 96692 40012
rect 96740 39956 96796 40012
rect 96844 39956 96900 40012
rect 127356 39956 127412 40012
rect 127460 39956 127516 40012
rect 127564 39956 127620 40012
rect 158076 39956 158132 40012
rect 158180 39956 158236 40012
rect 158284 39956 158340 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 81276 39172 81332 39228
rect 81380 39172 81436 39228
rect 81484 39172 81540 39228
rect 111996 39172 112052 39228
rect 112100 39172 112156 39228
rect 112204 39172 112260 39228
rect 142716 39172 142772 39228
rect 142820 39172 142876 39228
rect 142924 39172 142980 39228
rect 173436 39172 173492 39228
rect 173540 39172 173596 39228
rect 173644 39172 173700 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 96636 38388 96692 38444
rect 96740 38388 96796 38444
rect 96844 38388 96900 38444
rect 127356 38388 127412 38444
rect 127460 38388 127516 38444
rect 127564 38388 127620 38444
rect 158076 38388 158132 38444
rect 158180 38388 158236 38444
rect 158284 38388 158340 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 81276 37604 81332 37660
rect 81380 37604 81436 37660
rect 81484 37604 81540 37660
rect 111996 37604 112052 37660
rect 112100 37604 112156 37660
rect 112204 37604 112260 37660
rect 142716 37604 142772 37660
rect 142820 37604 142876 37660
rect 142924 37604 142980 37660
rect 173436 37604 173492 37660
rect 173540 37604 173596 37660
rect 173644 37604 173700 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 96636 36820 96692 36876
rect 96740 36820 96796 36876
rect 96844 36820 96900 36876
rect 127356 36820 127412 36876
rect 127460 36820 127516 36876
rect 127564 36820 127620 36876
rect 158076 36820 158132 36876
rect 158180 36820 158236 36876
rect 158284 36820 158340 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 81276 36036 81332 36092
rect 81380 36036 81436 36092
rect 81484 36036 81540 36092
rect 111996 36036 112052 36092
rect 112100 36036 112156 36092
rect 112204 36036 112260 36092
rect 142716 36036 142772 36092
rect 142820 36036 142876 36092
rect 142924 36036 142980 36092
rect 173436 36036 173492 36092
rect 173540 36036 173596 36092
rect 173644 36036 173700 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 96636 35252 96692 35308
rect 96740 35252 96796 35308
rect 96844 35252 96900 35308
rect 127356 35252 127412 35308
rect 127460 35252 127516 35308
rect 127564 35252 127620 35308
rect 158076 35252 158132 35308
rect 158180 35252 158236 35308
rect 158284 35252 158340 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 81276 34468 81332 34524
rect 81380 34468 81436 34524
rect 81484 34468 81540 34524
rect 111996 34468 112052 34524
rect 112100 34468 112156 34524
rect 112204 34468 112260 34524
rect 142716 34468 142772 34524
rect 142820 34468 142876 34524
rect 142924 34468 142980 34524
rect 173436 34468 173492 34524
rect 173540 34468 173596 34524
rect 173644 34468 173700 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 96636 33684 96692 33740
rect 96740 33684 96796 33740
rect 96844 33684 96900 33740
rect 127356 33684 127412 33740
rect 127460 33684 127516 33740
rect 127564 33684 127620 33740
rect 158076 33684 158132 33740
rect 158180 33684 158236 33740
rect 158284 33684 158340 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 81276 32900 81332 32956
rect 81380 32900 81436 32956
rect 81484 32900 81540 32956
rect 111996 32900 112052 32956
rect 112100 32900 112156 32956
rect 112204 32900 112260 32956
rect 142716 32900 142772 32956
rect 142820 32900 142876 32956
rect 142924 32900 142980 32956
rect 173436 32900 173492 32956
rect 173540 32900 173596 32956
rect 173644 32900 173700 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 96636 32116 96692 32172
rect 96740 32116 96796 32172
rect 96844 32116 96900 32172
rect 127356 32116 127412 32172
rect 127460 32116 127516 32172
rect 127564 32116 127620 32172
rect 158076 32116 158132 32172
rect 158180 32116 158236 32172
rect 158284 32116 158340 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 81276 31332 81332 31388
rect 81380 31332 81436 31388
rect 81484 31332 81540 31388
rect 111996 31332 112052 31388
rect 112100 31332 112156 31388
rect 112204 31332 112260 31388
rect 142716 31332 142772 31388
rect 142820 31332 142876 31388
rect 142924 31332 142980 31388
rect 173436 31332 173492 31388
rect 173540 31332 173596 31388
rect 173644 31332 173700 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 96636 30548 96692 30604
rect 96740 30548 96796 30604
rect 96844 30548 96900 30604
rect 127356 30548 127412 30604
rect 127460 30548 127516 30604
rect 127564 30548 127620 30604
rect 158076 30548 158132 30604
rect 158180 30548 158236 30604
rect 158284 30548 158340 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 81276 29764 81332 29820
rect 81380 29764 81436 29820
rect 81484 29764 81540 29820
rect 111996 29764 112052 29820
rect 112100 29764 112156 29820
rect 112204 29764 112260 29820
rect 142716 29764 142772 29820
rect 142820 29764 142876 29820
rect 142924 29764 142980 29820
rect 173436 29764 173492 29820
rect 173540 29764 173596 29820
rect 173644 29764 173700 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 96636 28980 96692 29036
rect 96740 28980 96796 29036
rect 96844 28980 96900 29036
rect 127356 28980 127412 29036
rect 127460 28980 127516 29036
rect 127564 28980 127620 29036
rect 158076 28980 158132 29036
rect 158180 28980 158236 29036
rect 158284 28980 158340 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 81276 28196 81332 28252
rect 81380 28196 81436 28252
rect 81484 28196 81540 28252
rect 111996 28196 112052 28252
rect 112100 28196 112156 28252
rect 112204 28196 112260 28252
rect 142716 28196 142772 28252
rect 142820 28196 142876 28252
rect 142924 28196 142980 28252
rect 173436 28196 173492 28252
rect 173540 28196 173596 28252
rect 173644 28196 173700 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 96636 27412 96692 27468
rect 96740 27412 96796 27468
rect 96844 27412 96900 27468
rect 127356 27412 127412 27468
rect 127460 27412 127516 27468
rect 127564 27412 127620 27468
rect 158076 27412 158132 27468
rect 158180 27412 158236 27468
rect 158284 27412 158340 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 81276 26628 81332 26684
rect 81380 26628 81436 26684
rect 81484 26628 81540 26684
rect 111996 26628 112052 26684
rect 112100 26628 112156 26684
rect 112204 26628 112260 26684
rect 142716 26628 142772 26684
rect 142820 26628 142876 26684
rect 142924 26628 142980 26684
rect 173436 26628 173492 26684
rect 173540 26628 173596 26684
rect 173644 26628 173700 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 96636 25844 96692 25900
rect 96740 25844 96796 25900
rect 96844 25844 96900 25900
rect 127356 25844 127412 25900
rect 127460 25844 127516 25900
rect 127564 25844 127620 25900
rect 158076 25844 158132 25900
rect 158180 25844 158236 25900
rect 158284 25844 158340 25900
rect 124236 25340 124292 25396
rect 127708 25228 127764 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 81276 25060 81332 25116
rect 81380 25060 81436 25116
rect 81484 25060 81540 25116
rect 111996 25060 112052 25116
rect 112100 25060 112156 25116
rect 112204 25060 112260 25116
rect 142716 25060 142772 25116
rect 142820 25060 142876 25116
rect 142924 25060 142980 25116
rect 173436 25060 173492 25116
rect 173540 25060 173596 25116
rect 173644 25060 173700 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 96636 24276 96692 24332
rect 96740 24276 96796 24332
rect 96844 24276 96900 24332
rect 127356 24276 127412 24332
rect 127460 24276 127516 24332
rect 127564 24276 127620 24332
rect 158076 24276 158132 24332
rect 158180 24276 158236 24332
rect 158284 24276 158340 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 81276 23492 81332 23548
rect 81380 23492 81436 23548
rect 81484 23492 81540 23548
rect 111996 23492 112052 23548
rect 112100 23492 112156 23548
rect 112204 23492 112260 23548
rect 142716 23492 142772 23548
rect 142820 23492 142876 23548
rect 142924 23492 142980 23548
rect 173436 23492 173492 23548
rect 173540 23492 173596 23548
rect 173644 23492 173700 23548
rect 113148 22876 113204 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 96636 22708 96692 22764
rect 96740 22708 96796 22764
rect 96844 22708 96900 22764
rect 127356 22708 127412 22764
rect 127460 22708 127516 22764
rect 127564 22708 127620 22764
rect 158076 22708 158132 22764
rect 158180 22708 158236 22764
rect 158284 22708 158340 22764
rect 83916 22652 83972 22708
rect 84476 22540 84532 22596
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 81276 21924 81332 21980
rect 81380 21924 81436 21980
rect 81484 21924 81540 21980
rect 111996 21924 112052 21980
rect 112100 21924 112156 21980
rect 112204 21924 112260 21980
rect 142716 21924 142772 21980
rect 142820 21924 142876 21980
rect 142924 21924 142980 21980
rect 173436 21924 173492 21980
rect 173540 21924 173596 21980
rect 173644 21924 173700 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 96636 21140 96692 21196
rect 96740 21140 96796 21196
rect 96844 21140 96900 21196
rect 127356 21140 127412 21196
rect 127460 21140 127516 21196
rect 127564 21140 127620 21196
rect 158076 21140 158132 21196
rect 158180 21140 158236 21196
rect 158284 21140 158340 21196
rect 123676 20524 123732 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 81276 20356 81332 20412
rect 81380 20356 81436 20412
rect 81484 20356 81540 20412
rect 111996 20356 112052 20412
rect 112100 20356 112156 20412
rect 112204 20356 112260 20412
rect 142716 20356 142772 20412
rect 142820 20356 142876 20412
rect 142924 20356 142980 20412
rect 173436 20356 173492 20412
rect 173540 20356 173596 20412
rect 173644 20356 173700 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 96636 19572 96692 19628
rect 96740 19572 96796 19628
rect 96844 19572 96900 19628
rect 127356 19572 127412 19628
rect 127460 19572 127516 19628
rect 127564 19572 127620 19628
rect 158076 19572 158132 19628
rect 158180 19572 158236 19628
rect 158284 19572 158340 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 81276 18788 81332 18844
rect 81380 18788 81436 18844
rect 81484 18788 81540 18844
rect 111996 18788 112052 18844
rect 112100 18788 112156 18844
rect 112204 18788 112260 18844
rect 142716 18788 142772 18844
rect 142820 18788 142876 18844
rect 142924 18788 142980 18844
rect 173436 18788 173492 18844
rect 173540 18788 173596 18844
rect 173644 18788 173700 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 96636 18004 96692 18060
rect 96740 18004 96796 18060
rect 96844 18004 96900 18060
rect 127356 18004 127412 18060
rect 127460 18004 127516 18060
rect 127564 18004 127620 18060
rect 158076 18004 158132 18060
rect 158180 18004 158236 18060
rect 158284 18004 158340 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 81276 17220 81332 17276
rect 81380 17220 81436 17276
rect 81484 17220 81540 17276
rect 111996 17220 112052 17276
rect 112100 17220 112156 17276
rect 112204 17220 112260 17276
rect 142716 17220 142772 17276
rect 142820 17220 142876 17276
rect 142924 17220 142980 17276
rect 173436 17220 173492 17276
rect 173540 17220 173596 17276
rect 173644 17220 173700 17276
rect 121212 16940 121268 16996
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 96636 16436 96692 16492
rect 96740 16436 96796 16492
rect 96844 16436 96900 16492
rect 127356 16436 127412 16492
rect 127460 16436 127516 16492
rect 127564 16436 127620 16492
rect 158076 16436 158132 16492
rect 158180 16436 158236 16492
rect 158284 16436 158340 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 81276 15652 81332 15708
rect 81380 15652 81436 15708
rect 81484 15652 81540 15708
rect 111996 15652 112052 15708
rect 112100 15652 112156 15708
rect 112204 15652 112260 15708
rect 142716 15652 142772 15708
rect 142820 15652 142876 15708
rect 142924 15652 142980 15708
rect 173436 15652 173492 15708
rect 173540 15652 173596 15708
rect 173644 15652 173700 15708
rect 128156 15260 128212 15316
rect 85596 15148 85652 15204
rect 137004 15148 137060 15204
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 96636 14868 96692 14924
rect 96740 14868 96796 14924
rect 96844 14868 96900 14924
rect 127356 14868 127412 14924
rect 127460 14868 127516 14924
rect 127564 14868 127620 14924
rect 158076 14868 158132 14924
rect 158180 14868 158236 14924
rect 158284 14868 158340 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 81276 14084 81332 14140
rect 81380 14084 81436 14140
rect 81484 14084 81540 14140
rect 111996 14084 112052 14140
rect 112100 14084 112156 14140
rect 112204 14084 112260 14140
rect 142716 14084 142772 14140
rect 142820 14084 142876 14140
rect 142924 14084 142980 14140
rect 173436 14084 173492 14140
rect 173540 14084 173596 14140
rect 173644 14084 173700 14140
rect 111804 14028 111860 14084
rect 79884 13692 79940 13748
rect 68348 13580 68404 13636
rect 77420 13580 77476 13636
rect 78652 13580 78708 13636
rect 91532 13692 91588 13748
rect 111804 13580 111860 13636
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 96636 13300 96692 13356
rect 96740 13300 96796 13356
rect 96844 13300 96900 13356
rect 127356 13300 127412 13356
rect 127460 13300 127516 13356
rect 127564 13300 127620 13356
rect 158076 13300 158132 13356
rect 158180 13300 158236 13356
rect 158284 13300 158340 13356
rect 69356 13020 69412 13076
rect 74732 12684 74788 12740
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 81276 12516 81332 12572
rect 81380 12516 81436 12572
rect 81484 12516 81540 12572
rect 111996 12516 112052 12572
rect 112100 12516 112156 12572
rect 112204 12516 112260 12572
rect 142716 12516 142772 12572
rect 142820 12516 142876 12572
rect 142924 12516 142980 12572
rect 173436 12516 173492 12572
rect 173540 12516 173596 12572
rect 173644 12516 173700 12572
rect 70252 12348 70308 12404
rect 83356 12012 83412 12068
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 96636 11732 96692 11788
rect 96740 11732 96796 11788
rect 96844 11732 96900 11788
rect 127356 11732 127412 11788
rect 127460 11732 127516 11788
rect 127564 11732 127620 11788
rect 158076 11732 158132 11788
rect 158180 11732 158236 11788
rect 158284 11732 158340 11788
rect 97020 11564 97076 11620
rect 63756 11452 63812 11508
rect 99820 11116 99876 11172
rect 113260 11116 113316 11172
rect 114716 11116 114772 11172
rect 99484 11004 99540 11060
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 81276 10948 81332 11004
rect 81380 10948 81436 11004
rect 81484 10948 81540 11004
rect 111996 10948 112052 11004
rect 112100 10948 112156 11004
rect 112204 10948 112260 11004
rect 142716 10948 142772 11004
rect 142820 10948 142876 11004
rect 142924 10948 142980 11004
rect 173436 10948 173492 11004
rect 173540 10948 173596 11004
rect 173644 10948 173700 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 99708 10444 99764 10500
rect 117292 10444 117348 10500
rect 99484 10332 99540 10388
rect 109788 10332 109844 10388
rect 97020 10220 97076 10276
rect 99596 10220 99652 10276
rect 109340 10220 109396 10276
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 96636 10164 96692 10220
rect 96740 10164 96796 10220
rect 96844 10164 96900 10220
rect 127356 10164 127412 10220
rect 127460 10164 127516 10220
rect 127564 10164 127620 10220
rect 158076 10164 158132 10220
rect 158180 10164 158236 10220
rect 158284 10164 158340 10220
rect 114492 10108 114548 10164
rect 135660 10108 135716 10164
rect 96348 9996 96404 10052
rect 106764 9996 106820 10052
rect 84476 9884 84532 9940
rect 113932 9772 113988 9828
rect 119756 9772 119812 9828
rect 104188 9548 104244 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 81276 9380 81332 9436
rect 81380 9380 81436 9436
rect 81484 9380 81540 9436
rect 111996 9380 112052 9436
rect 112100 9380 112156 9436
rect 112204 9380 112260 9436
rect 142716 9380 142772 9436
rect 142820 9380 142876 9436
rect 142924 9380 142980 9436
rect 173436 9380 173492 9436
rect 173540 9380 173596 9436
rect 173644 9380 173700 9436
rect 94444 9212 94500 9268
rect 121212 9212 121268 9268
rect 78316 8652 78372 8708
rect 102172 8652 102228 8708
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 96636 8596 96692 8652
rect 96740 8596 96796 8652
rect 96844 8596 96900 8652
rect 127356 8596 127412 8652
rect 127460 8596 127516 8652
rect 127564 8596 127620 8652
rect 158076 8596 158132 8652
rect 158180 8596 158236 8652
rect 158284 8596 158340 8652
rect 95676 8428 95732 8484
rect 102396 8316 102452 8372
rect 136668 8204 136724 8260
rect 77868 7980 77924 8036
rect 102396 7980 102452 8036
rect 62300 7868 62356 7924
rect 63756 7868 63812 7924
rect 96124 7868 96180 7924
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 81276 7812 81332 7868
rect 81380 7812 81436 7868
rect 81484 7812 81540 7868
rect 111996 7812 112052 7868
rect 112100 7812 112156 7868
rect 112204 7812 112260 7868
rect 142716 7812 142772 7868
rect 142820 7812 142876 7868
rect 142924 7812 142980 7868
rect 173436 7812 173492 7868
rect 173540 7812 173596 7868
rect 173644 7812 173700 7868
rect 94444 7644 94500 7700
rect 121324 7644 121380 7700
rect 67116 7532 67172 7588
rect 95676 7532 95732 7588
rect 77868 7308 77924 7364
rect 83916 7308 83972 7364
rect 96124 7308 96180 7364
rect 140476 7308 140532 7364
rect 113932 7196 113988 7252
rect 114716 7196 114772 7252
rect 82124 7084 82180 7140
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 96636 7028 96692 7084
rect 96740 7028 96796 7084
rect 96844 7028 96900 7084
rect 127356 7028 127412 7084
rect 127460 7028 127516 7084
rect 127564 7028 127620 7084
rect 158076 7028 158132 7084
rect 158180 7028 158236 7084
rect 158284 7028 158340 7084
rect 137340 6972 137396 7028
rect 122108 6748 122164 6804
rect 137564 6748 137620 6804
rect 57148 6636 57204 6692
rect 84476 6636 84532 6692
rect 91532 6636 91588 6692
rect 104188 6636 104244 6692
rect 106764 6636 106820 6692
rect 78316 6524 78372 6580
rect 136668 6524 136724 6580
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 79884 6300 79940 6356
rect 82124 6300 82180 6356
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 81276 6244 81332 6300
rect 81380 6244 81436 6300
rect 81484 6244 81540 6300
rect 111996 6244 112052 6300
rect 112100 6244 112156 6300
rect 112204 6244 112260 6300
rect 116396 6188 116452 6244
rect 142716 6244 142772 6300
rect 142820 6244 142876 6300
rect 142924 6244 142980 6300
rect 173436 6244 173492 6300
rect 173540 6244 173596 6300
rect 173644 6244 173700 6300
rect 132972 6188 133028 6244
rect 137340 6188 137396 6244
rect 137004 6076 137060 6132
rect 69356 5964 69412 6020
rect 123676 5964 123732 6020
rect 134652 5852 134708 5908
rect 74732 5740 74788 5796
rect 116396 5740 116452 5796
rect 136668 5740 136724 5796
rect 79884 5628 79940 5684
rect 102396 5628 102452 5684
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 96636 5460 96692 5516
rect 96740 5460 96796 5516
rect 96844 5460 96900 5516
rect 135660 5628 135716 5684
rect 127356 5460 127412 5516
rect 127460 5460 127516 5516
rect 127564 5460 127620 5516
rect 133868 5404 133924 5460
rect 135884 5404 135940 5460
rect 158076 5460 158132 5516
rect 158180 5460 158236 5516
rect 158284 5460 158340 5516
rect 78652 5180 78708 5236
rect 95340 5180 95396 5236
rect 99820 5180 99876 5236
rect 70252 5068 70308 5124
rect 96348 5068 96404 5124
rect 119756 5068 119812 5124
rect 111804 4956 111860 5012
rect 122108 4956 122164 5012
rect 69132 4732 69188 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 81276 4676 81332 4732
rect 81380 4676 81436 4732
rect 81484 4676 81540 4732
rect 83356 4844 83412 4900
rect 91420 4844 91476 4900
rect 111804 4732 111860 4788
rect 113932 4732 113988 4788
rect 111996 4676 112052 4732
rect 112100 4676 112156 4732
rect 112204 4676 112260 4732
rect 142716 4676 142772 4732
rect 142820 4676 142876 4732
rect 142924 4676 142980 4732
rect 62300 4620 62356 4676
rect 77420 4620 77476 4676
rect 91308 4620 91364 4676
rect 67116 4396 67172 4452
rect 68348 4396 68404 4452
rect 69132 4396 69188 4452
rect 113260 4508 113316 4564
rect 117292 4508 117348 4564
rect 127708 4508 127764 4564
rect 135660 4508 135716 4564
rect 135884 4508 135940 4564
rect 104188 4396 104244 4452
rect 85596 4284 85652 4340
rect 102172 4284 102228 4340
rect 173436 4676 173492 4732
rect 173540 4676 173596 4732
rect 173644 4676 173700 4732
rect 121324 4284 121380 4340
rect 114492 4172 114548 4228
rect 133868 4172 133924 4228
rect 134652 4172 134708 4228
rect 140476 4060 140532 4116
rect 137564 3948 137620 4004
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 96636 3892 96692 3948
rect 96740 3892 96796 3948
rect 96844 3892 96900 3948
rect 127356 3892 127412 3948
rect 127460 3892 127516 3948
rect 127564 3892 127620 3948
rect 158076 3892 158132 3948
rect 158180 3892 158236 3948
rect 158284 3892 158340 3948
rect 121772 3836 121828 3892
rect 121548 3724 121604 3780
rect 132972 3724 133028 3780
rect 121212 3500 121268 3556
rect 124236 3276 124292 3332
rect 128156 3276 128212 3332
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 81276 3108 81332 3164
rect 81380 3108 81436 3164
rect 81484 3108 81540 3164
rect 111996 3108 112052 3164
rect 112100 3108 112156 3164
rect 112204 3108 112260 3164
rect 142716 3108 142772 3164
rect 142820 3108 142876 3164
rect 142924 3108 142980 3164
rect 173436 3108 173492 3164
rect 173540 3108 173596 3164
rect 173644 3108 173700 3164
rect 117292 2940 117348 2996
<< metal4 >>
rect 4448 116844 4768 116876
rect 4448 116788 4476 116844
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4740 116788 4768 116844
rect 4448 115276 4768 116788
rect 4448 115220 4476 115276
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4740 115220 4768 115276
rect 4448 113708 4768 115220
rect 4448 113652 4476 113708
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4740 113652 4768 113708
rect 4448 112140 4768 113652
rect 4448 112084 4476 112140
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4740 112084 4768 112140
rect 4448 110572 4768 112084
rect 4448 110516 4476 110572
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4740 110516 4768 110572
rect 4448 109004 4768 110516
rect 4448 108948 4476 109004
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4740 108948 4768 109004
rect 4448 107436 4768 108948
rect 4448 107380 4476 107436
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4740 107380 4768 107436
rect 4448 105868 4768 107380
rect 4448 105812 4476 105868
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4740 105812 4768 105868
rect 4448 104300 4768 105812
rect 4448 104244 4476 104300
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4740 104244 4768 104300
rect 4448 102732 4768 104244
rect 4448 102676 4476 102732
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4740 102676 4768 102732
rect 4448 101164 4768 102676
rect 4448 101108 4476 101164
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4740 101108 4768 101164
rect 4448 99596 4768 101108
rect 4448 99540 4476 99596
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4740 99540 4768 99596
rect 4448 98028 4768 99540
rect 4448 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4768 98028
rect 4448 96460 4768 97972
rect 4448 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4768 96460
rect 4448 94892 4768 96404
rect 4448 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4768 94892
rect 4448 93324 4768 94836
rect 4448 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4768 93324
rect 4448 91756 4768 93268
rect 4448 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4768 91756
rect 4448 90188 4768 91700
rect 4448 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4768 90188
rect 4448 88620 4768 90132
rect 4448 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4768 88620
rect 4448 87052 4768 88564
rect 4448 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4768 87052
rect 4448 85484 4768 86996
rect 4448 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4768 85484
rect 4448 83916 4768 85428
rect 4448 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4768 83916
rect 4448 82348 4768 83860
rect 4448 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4768 82348
rect 4448 80780 4768 82292
rect 4448 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4768 80780
rect 4448 79212 4768 80724
rect 4448 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4768 79212
rect 4448 77644 4768 79156
rect 4448 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4768 77644
rect 4448 76076 4768 77588
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 116060 20128 116876
rect 19808 116004 19836 116060
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 20100 116004 20128 116060
rect 19808 114492 20128 116004
rect 19808 114436 19836 114492
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 20100 114436 20128 114492
rect 19808 112924 20128 114436
rect 19808 112868 19836 112924
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 20100 112868 20128 112924
rect 19808 111356 20128 112868
rect 19808 111300 19836 111356
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 20100 111300 20128 111356
rect 19808 109788 20128 111300
rect 19808 109732 19836 109788
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 20100 109732 20128 109788
rect 19808 108220 20128 109732
rect 19808 108164 19836 108220
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 20100 108164 20128 108220
rect 19808 106652 20128 108164
rect 19808 106596 19836 106652
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 20100 106596 20128 106652
rect 19808 105084 20128 106596
rect 19808 105028 19836 105084
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 20100 105028 20128 105084
rect 19808 103516 20128 105028
rect 19808 103460 19836 103516
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 20100 103460 20128 103516
rect 19808 101948 20128 103460
rect 19808 101892 19836 101948
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 20100 101892 20128 101948
rect 19808 100380 20128 101892
rect 19808 100324 19836 100380
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 20100 100324 20128 100380
rect 19808 98812 20128 100324
rect 19808 98756 19836 98812
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 20100 98756 20128 98812
rect 19808 97244 20128 98756
rect 19808 97188 19836 97244
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 20100 97188 20128 97244
rect 19808 95676 20128 97188
rect 19808 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20128 95676
rect 19808 94108 20128 95620
rect 19808 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20128 94108
rect 19808 92540 20128 94052
rect 19808 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20128 92540
rect 19808 90972 20128 92484
rect 19808 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20128 90972
rect 19808 89404 20128 90916
rect 19808 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20128 89404
rect 19808 87836 20128 89348
rect 19808 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20128 87836
rect 19808 86268 20128 87780
rect 19808 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20128 86268
rect 19808 84700 20128 86212
rect 19808 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20128 84700
rect 19808 83132 20128 84644
rect 19808 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20128 83132
rect 19808 81564 20128 83076
rect 19808 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20128 81564
rect 19808 79996 20128 81508
rect 19808 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20128 79996
rect 19808 78428 20128 79940
rect 19808 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20128 78428
rect 19808 76860 20128 78372
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 116844 35488 116876
rect 35168 116788 35196 116844
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35460 116788 35488 116844
rect 35168 115276 35488 116788
rect 35168 115220 35196 115276
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35460 115220 35488 115276
rect 35168 113708 35488 115220
rect 35168 113652 35196 113708
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35460 113652 35488 113708
rect 35168 112140 35488 113652
rect 35168 112084 35196 112140
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35460 112084 35488 112140
rect 35168 110572 35488 112084
rect 35168 110516 35196 110572
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35460 110516 35488 110572
rect 35168 109004 35488 110516
rect 35168 108948 35196 109004
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35460 108948 35488 109004
rect 35168 107436 35488 108948
rect 35168 107380 35196 107436
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35460 107380 35488 107436
rect 35168 105868 35488 107380
rect 35168 105812 35196 105868
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35460 105812 35488 105868
rect 35168 104300 35488 105812
rect 35168 104244 35196 104300
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35460 104244 35488 104300
rect 35168 102732 35488 104244
rect 35168 102676 35196 102732
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35460 102676 35488 102732
rect 35168 101164 35488 102676
rect 35168 101108 35196 101164
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35460 101108 35488 101164
rect 35168 99596 35488 101108
rect 35168 99540 35196 99596
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35460 99540 35488 99596
rect 35168 98028 35488 99540
rect 35168 97972 35196 98028
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35460 97972 35488 98028
rect 35168 96460 35488 97972
rect 35168 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35488 96460
rect 35168 94892 35488 96404
rect 35168 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35488 94892
rect 35168 93324 35488 94836
rect 35168 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35488 93324
rect 35168 91756 35488 93268
rect 35168 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35488 91756
rect 35168 90188 35488 91700
rect 35168 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35488 90188
rect 35168 88620 35488 90132
rect 35168 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35488 88620
rect 35168 87052 35488 88564
rect 35168 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35488 87052
rect 35168 85484 35488 86996
rect 35168 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35488 85484
rect 35168 83916 35488 85428
rect 35168 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35488 83916
rect 35168 82348 35488 83860
rect 35168 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35488 82348
rect 35168 80780 35488 82292
rect 35168 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35488 80780
rect 35168 79212 35488 80724
rect 35168 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35488 79212
rect 35168 77644 35488 79156
rect 35168 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35488 77644
rect 35168 76076 35488 77588
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 116060 50848 116876
rect 50528 116004 50556 116060
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50820 116004 50848 116060
rect 50528 114492 50848 116004
rect 50528 114436 50556 114492
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50820 114436 50848 114492
rect 50528 112924 50848 114436
rect 50528 112868 50556 112924
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50820 112868 50848 112924
rect 50528 111356 50848 112868
rect 50528 111300 50556 111356
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50820 111300 50848 111356
rect 50528 109788 50848 111300
rect 50528 109732 50556 109788
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50820 109732 50848 109788
rect 50528 108220 50848 109732
rect 65888 116844 66208 116876
rect 65888 116788 65916 116844
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 66180 116788 66208 116844
rect 65888 115276 66208 116788
rect 65888 115220 65916 115276
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 66180 115220 66208 115276
rect 65888 113708 66208 115220
rect 65888 113652 65916 113708
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 66180 113652 66208 113708
rect 65888 112140 66208 113652
rect 65888 112084 65916 112140
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 66180 112084 66208 112140
rect 65888 110572 66208 112084
rect 65888 110516 65916 110572
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 66180 110516 66208 110572
rect 65888 109004 66208 110516
rect 65888 108948 65916 109004
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 66180 108948 66208 109004
rect 50528 108164 50556 108220
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50820 108164 50848 108220
rect 50528 106652 50848 108164
rect 50528 106596 50556 106652
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50820 106596 50848 106652
rect 50528 105084 50848 106596
rect 50528 105028 50556 105084
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50820 105028 50848 105084
rect 50528 103516 50848 105028
rect 50528 103460 50556 103516
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50820 103460 50848 103516
rect 50528 101948 50848 103460
rect 50528 101892 50556 101948
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50820 101892 50848 101948
rect 50528 100380 50848 101892
rect 50528 100324 50556 100380
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50820 100324 50848 100380
rect 50528 98812 50848 100324
rect 50528 98756 50556 98812
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50820 98756 50848 98812
rect 50528 97244 50848 98756
rect 50528 97188 50556 97244
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50820 97188 50848 97244
rect 50528 95676 50848 97188
rect 50528 95620 50556 95676
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50820 95620 50848 95676
rect 50528 94108 50848 95620
rect 50528 94052 50556 94108
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50820 94052 50848 94108
rect 50528 92540 50848 94052
rect 50528 92484 50556 92540
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50820 92484 50848 92540
rect 50528 90972 50848 92484
rect 50528 90916 50556 90972
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50820 90916 50848 90972
rect 50528 89404 50848 90916
rect 50528 89348 50556 89404
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50820 89348 50848 89404
rect 50528 87836 50848 89348
rect 50528 87780 50556 87836
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50820 87780 50848 87836
rect 50528 86268 50848 87780
rect 50528 86212 50556 86268
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50820 86212 50848 86268
rect 50528 84700 50848 86212
rect 50528 84644 50556 84700
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50820 84644 50848 84700
rect 50528 83132 50848 84644
rect 50528 83076 50556 83132
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50820 83076 50848 83132
rect 50528 81564 50848 83076
rect 50528 81508 50556 81564
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50820 81508 50848 81564
rect 50528 79996 50848 81508
rect 50528 79940 50556 79996
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50820 79940 50848 79996
rect 50528 78428 50848 79940
rect 50528 78372 50556 78428
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50820 78372 50848 78428
rect 50528 76860 50848 78372
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 57148 108388 57204 108398
rect 57148 6692 57204 108332
rect 65888 107436 66208 108948
rect 65888 107380 65916 107436
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 66180 107380 66208 107436
rect 65888 105868 66208 107380
rect 65888 105812 65916 105868
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 66180 105812 66208 105868
rect 65888 104300 66208 105812
rect 65888 104244 65916 104300
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 66180 104244 66208 104300
rect 65888 102732 66208 104244
rect 65888 102676 65916 102732
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 66180 102676 66208 102732
rect 65888 101164 66208 102676
rect 65888 101108 65916 101164
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 66180 101108 66208 101164
rect 65888 99596 66208 101108
rect 65888 99540 65916 99596
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 66180 99540 66208 99596
rect 65888 98028 66208 99540
rect 65888 97972 65916 98028
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 66180 97972 66208 98028
rect 65888 96460 66208 97972
rect 65888 96404 65916 96460
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 66180 96404 66208 96460
rect 65888 94892 66208 96404
rect 65888 94836 65916 94892
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 66180 94836 66208 94892
rect 65888 93324 66208 94836
rect 65888 93268 65916 93324
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 66180 93268 66208 93324
rect 65888 91756 66208 93268
rect 65888 91700 65916 91756
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 66180 91700 66208 91756
rect 65888 90188 66208 91700
rect 65888 90132 65916 90188
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 66180 90132 66208 90188
rect 65888 88620 66208 90132
rect 65888 88564 65916 88620
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 66180 88564 66208 88620
rect 65888 87052 66208 88564
rect 65888 86996 65916 87052
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 66180 86996 66208 87052
rect 65888 85484 66208 86996
rect 65888 85428 65916 85484
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 66180 85428 66208 85484
rect 65888 83916 66208 85428
rect 65888 83860 65916 83916
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 66180 83860 66208 83916
rect 65888 82348 66208 83860
rect 65888 82292 65916 82348
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 66180 82292 66208 82348
rect 65888 80780 66208 82292
rect 65888 80724 65916 80780
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 66180 80724 66208 80780
rect 65888 79212 66208 80724
rect 65888 79156 65916 79212
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 66180 79156 66208 79212
rect 65888 77644 66208 79156
rect 65888 77588 65916 77644
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 66180 77588 66208 77644
rect 65888 76076 66208 77588
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 81248 116060 81568 116876
rect 96608 116844 96928 116876
rect 96608 116788 96636 116844
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96900 116788 96928 116844
rect 81248 116004 81276 116060
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81540 116004 81568 116060
rect 81248 114492 81568 116004
rect 81248 114436 81276 114492
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81540 114436 81568 114492
rect 81248 112924 81568 114436
rect 81248 112868 81276 112924
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81540 112868 81568 112924
rect 81248 111356 81568 112868
rect 81248 111300 81276 111356
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81540 111300 81568 111356
rect 81248 109788 81568 111300
rect 81248 109732 81276 109788
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81540 109732 81568 109788
rect 81248 108220 81568 109732
rect 81248 108164 81276 108220
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81540 108164 81568 108220
rect 81248 106652 81568 108164
rect 81248 106596 81276 106652
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81540 106596 81568 106652
rect 81248 105084 81568 106596
rect 81248 105028 81276 105084
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81540 105028 81568 105084
rect 81248 103516 81568 105028
rect 81248 103460 81276 103516
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81540 103460 81568 103516
rect 81248 101948 81568 103460
rect 81248 101892 81276 101948
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81540 101892 81568 101948
rect 81248 100380 81568 101892
rect 81248 100324 81276 100380
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81540 100324 81568 100380
rect 81248 98812 81568 100324
rect 81248 98756 81276 98812
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81540 98756 81568 98812
rect 81248 97244 81568 98756
rect 81248 97188 81276 97244
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81540 97188 81568 97244
rect 81248 95676 81568 97188
rect 81248 95620 81276 95676
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81540 95620 81568 95676
rect 81248 94108 81568 95620
rect 81248 94052 81276 94108
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81540 94052 81568 94108
rect 81248 92540 81568 94052
rect 81248 92484 81276 92540
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81540 92484 81568 92540
rect 81248 90972 81568 92484
rect 81248 90916 81276 90972
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81540 90916 81568 90972
rect 81248 89404 81568 90916
rect 81248 89348 81276 89404
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81540 89348 81568 89404
rect 81248 87836 81568 89348
rect 81248 87780 81276 87836
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81540 87780 81568 87836
rect 81248 86268 81568 87780
rect 81248 86212 81276 86268
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81540 86212 81568 86268
rect 81248 84700 81568 86212
rect 81248 84644 81276 84700
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81540 84644 81568 84700
rect 81248 83132 81568 84644
rect 81248 83076 81276 83132
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81540 83076 81568 83132
rect 81248 81564 81568 83076
rect 81248 81508 81276 81564
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81540 81508 81568 81564
rect 81248 79996 81568 81508
rect 81248 79940 81276 79996
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81540 79940 81568 79996
rect 81248 78428 81568 79940
rect 81248 78372 81276 78428
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81540 78372 81568 78428
rect 81248 76860 81568 78372
rect 81248 76804 81276 76860
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81540 76804 81568 76860
rect 81248 75292 81568 76804
rect 81248 75236 81276 75292
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81540 75236 81568 75292
rect 81248 73724 81568 75236
rect 81248 73668 81276 73724
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81540 73668 81568 73724
rect 81248 72156 81568 73668
rect 81248 72100 81276 72156
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81540 72100 81568 72156
rect 81248 70588 81568 72100
rect 81248 70532 81276 70588
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81540 70532 81568 70588
rect 81248 69020 81568 70532
rect 81248 68964 81276 69020
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81540 68964 81568 69020
rect 81248 67452 81568 68964
rect 81248 67396 81276 67452
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81540 67396 81568 67452
rect 81248 65884 81568 67396
rect 81248 65828 81276 65884
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81540 65828 81568 65884
rect 81248 64316 81568 65828
rect 81248 64260 81276 64316
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81540 64260 81568 64316
rect 81248 62748 81568 64260
rect 81248 62692 81276 62748
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81540 62692 81568 62748
rect 81248 61180 81568 62692
rect 81248 61124 81276 61180
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81540 61124 81568 61180
rect 81248 59612 81568 61124
rect 81248 59556 81276 59612
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81540 59556 81568 59612
rect 81248 58044 81568 59556
rect 81248 57988 81276 58044
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81540 57988 81568 58044
rect 81248 56476 81568 57988
rect 81248 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81568 56476
rect 81248 54908 81568 56420
rect 81248 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81568 54908
rect 81248 53340 81568 54852
rect 81248 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81568 53340
rect 81248 51772 81568 53284
rect 81248 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81568 51772
rect 81248 50204 81568 51716
rect 81248 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81568 50204
rect 81248 48636 81568 50148
rect 81248 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81568 48636
rect 81248 47068 81568 48580
rect 81248 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81568 47068
rect 81248 45500 81568 47012
rect 81248 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81568 45500
rect 81248 43932 81568 45444
rect 81248 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81568 43932
rect 81248 42364 81568 43876
rect 81248 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81568 42364
rect 81248 40796 81568 42308
rect 81248 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81568 40796
rect 81248 39228 81568 40740
rect 81248 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81568 39228
rect 81248 37660 81568 39172
rect 81248 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81568 37660
rect 81248 36092 81568 37604
rect 81248 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81568 36092
rect 81248 34524 81568 36036
rect 81248 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81568 34524
rect 81248 32956 81568 34468
rect 81248 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81568 32956
rect 81248 31388 81568 32900
rect 81248 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81568 31388
rect 81248 29820 81568 31332
rect 81248 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81568 29820
rect 81248 28252 81568 29764
rect 81248 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81568 28252
rect 81248 26684 81568 28196
rect 81248 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81568 26684
rect 81248 25116 81568 26628
rect 81248 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81568 25116
rect 81248 23548 81568 25060
rect 81248 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81568 23548
rect 81248 21980 81568 23492
rect 95340 116228 95396 116238
rect 81248 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81568 21980
rect 81248 20412 81568 21924
rect 81248 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81568 20412
rect 81248 18844 81568 20356
rect 81248 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81568 18844
rect 81248 17276 81568 18788
rect 81248 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81568 17276
rect 81248 15708 81568 17220
rect 81248 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81568 15708
rect 81248 14140 81568 15652
rect 81248 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81568 14140
rect 79884 13748 79940 13758
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 63756 11508 63812 11518
rect 57148 6626 57204 6636
rect 62300 7924 62356 7934
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 62300 4676 62356 7868
rect 63756 7924 63812 11452
rect 63756 7858 63812 7868
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 62300 4610 62356 4620
rect 65888 7084 66208 8596
rect 68348 13636 68404 13646
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 3948 66208 5460
rect 67116 7588 67172 7598
rect 67116 4452 67172 7532
rect 67116 4386 67172 4396
rect 68348 4452 68404 13580
rect 77420 13636 77476 13646
rect 69356 13076 69412 13086
rect 69356 6020 69412 13020
rect 74732 12740 74788 12750
rect 69356 5954 69412 5964
rect 70252 12404 70308 12414
rect 70252 5124 70308 12348
rect 74732 5796 74788 12684
rect 74732 5730 74788 5740
rect 70252 5058 70308 5068
rect 68348 4386 68404 4396
rect 69132 4788 69188 4798
rect 69132 4452 69188 4732
rect 77420 4676 77476 13580
rect 78652 13636 78708 13646
rect 78316 8708 78372 8718
rect 77868 8036 77924 8046
rect 77868 7364 77924 7980
rect 77868 7298 77924 7308
rect 78316 6580 78372 8652
rect 78316 6514 78372 6524
rect 78652 5236 78708 13580
rect 79884 6356 79940 13692
rect 79884 5684 79940 6300
rect 79884 5618 79940 5628
rect 81248 12572 81568 14084
rect 81248 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81568 12572
rect 81248 11004 81568 12516
rect 83916 22708 83972 22718
rect 81248 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81568 11004
rect 81248 9436 81568 10948
rect 81248 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81568 9436
rect 81248 7868 81568 9380
rect 81248 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81568 7868
rect 81248 6300 81568 7812
rect 83356 12068 83412 12078
rect 81248 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81568 6300
rect 82124 7140 82180 7150
rect 82124 6356 82180 7084
rect 82124 6290 82180 6300
rect 78652 5170 78708 5180
rect 77420 4610 77476 4620
rect 81248 4732 81568 6244
rect 83356 4900 83412 12012
rect 83916 7364 83972 22652
rect 83916 7298 83972 7308
rect 84476 22596 84532 22606
rect 84476 9940 84532 22540
rect 84476 6692 84532 9884
rect 84476 6626 84532 6636
rect 85596 15204 85652 15214
rect 83356 4834 83412 4844
rect 81248 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81568 4732
rect 69132 4386 69188 4396
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
rect 81248 3164 81568 4676
rect 85596 4340 85652 15148
rect 91532 13748 91588 13758
rect 91532 6692 91588 13692
rect 94444 9268 94500 9278
rect 94444 7700 94500 9212
rect 94444 7634 94500 7644
rect 91532 6626 91588 6636
rect 95340 5236 95396 116172
rect 96608 115276 96928 116788
rect 96608 115220 96636 115276
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96900 115220 96928 115276
rect 96608 113708 96928 115220
rect 96608 113652 96636 113708
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96900 113652 96928 113708
rect 96608 112140 96928 113652
rect 96608 112084 96636 112140
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96900 112084 96928 112140
rect 96608 110572 96928 112084
rect 96608 110516 96636 110572
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96900 110516 96928 110572
rect 96608 109004 96928 110516
rect 96608 108948 96636 109004
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96900 108948 96928 109004
rect 96608 107436 96928 108948
rect 96608 107380 96636 107436
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96900 107380 96928 107436
rect 96608 105868 96928 107380
rect 96608 105812 96636 105868
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96900 105812 96928 105868
rect 96608 104300 96928 105812
rect 96608 104244 96636 104300
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96900 104244 96928 104300
rect 96608 102732 96928 104244
rect 96608 102676 96636 102732
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96900 102676 96928 102732
rect 96608 101164 96928 102676
rect 96608 101108 96636 101164
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96900 101108 96928 101164
rect 96608 99596 96928 101108
rect 96608 99540 96636 99596
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96900 99540 96928 99596
rect 96608 98028 96928 99540
rect 96608 97972 96636 98028
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96900 97972 96928 98028
rect 96608 96460 96928 97972
rect 96608 96404 96636 96460
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96900 96404 96928 96460
rect 96608 94892 96928 96404
rect 96608 94836 96636 94892
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96900 94836 96928 94892
rect 96608 93324 96928 94836
rect 96608 93268 96636 93324
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96900 93268 96928 93324
rect 96608 91756 96928 93268
rect 96608 91700 96636 91756
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96900 91700 96928 91756
rect 96608 90188 96928 91700
rect 96608 90132 96636 90188
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96900 90132 96928 90188
rect 96608 88620 96928 90132
rect 96608 88564 96636 88620
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96900 88564 96928 88620
rect 96608 87052 96928 88564
rect 96608 86996 96636 87052
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96900 86996 96928 87052
rect 96608 85484 96928 86996
rect 96608 85428 96636 85484
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96900 85428 96928 85484
rect 96608 83916 96928 85428
rect 96608 83860 96636 83916
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96900 83860 96928 83916
rect 96608 82348 96928 83860
rect 96608 82292 96636 82348
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96900 82292 96928 82348
rect 96608 80780 96928 82292
rect 96608 80724 96636 80780
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96900 80724 96928 80780
rect 96608 79212 96928 80724
rect 96608 79156 96636 79212
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96900 79156 96928 79212
rect 96608 77644 96928 79156
rect 96608 77588 96636 77644
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96900 77588 96928 77644
rect 96608 76076 96928 77588
rect 96608 76020 96636 76076
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96900 76020 96928 76076
rect 96608 74508 96928 76020
rect 96608 74452 96636 74508
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96900 74452 96928 74508
rect 96608 72940 96928 74452
rect 96608 72884 96636 72940
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96900 72884 96928 72940
rect 96608 71372 96928 72884
rect 96608 71316 96636 71372
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96900 71316 96928 71372
rect 96608 69804 96928 71316
rect 96608 69748 96636 69804
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96900 69748 96928 69804
rect 96608 68236 96928 69748
rect 96608 68180 96636 68236
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96900 68180 96928 68236
rect 96608 66668 96928 68180
rect 96608 66612 96636 66668
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96900 66612 96928 66668
rect 96608 65100 96928 66612
rect 96608 65044 96636 65100
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96900 65044 96928 65100
rect 96608 63532 96928 65044
rect 96608 63476 96636 63532
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96900 63476 96928 63532
rect 96608 61964 96928 63476
rect 96608 61908 96636 61964
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96900 61908 96928 61964
rect 96608 60396 96928 61908
rect 96608 60340 96636 60396
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96900 60340 96928 60396
rect 96608 58828 96928 60340
rect 96608 58772 96636 58828
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96900 58772 96928 58828
rect 96608 57260 96928 58772
rect 96608 57204 96636 57260
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96900 57204 96928 57260
rect 96608 55692 96928 57204
rect 96608 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96928 55692
rect 96608 54124 96928 55636
rect 96608 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96928 54124
rect 96608 52556 96928 54068
rect 96608 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96928 52556
rect 96608 50988 96928 52500
rect 96608 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96928 50988
rect 96608 49420 96928 50932
rect 96608 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96928 49420
rect 96608 47852 96928 49364
rect 96608 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96928 47852
rect 96608 46284 96928 47796
rect 96608 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96928 46284
rect 96608 44716 96928 46228
rect 96608 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96928 44716
rect 96608 43148 96928 44660
rect 96608 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96928 43148
rect 96608 41580 96928 43092
rect 96608 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96928 41580
rect 96608 40012 96928 41524
rect 96608 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96928 40012
rect 96608 38444 96928 39956
rect 96608 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96928 38444
rect 96608 36876 96928 38388
rect 96608 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96928 36876
rect 96608 35308 96928 36820
rect 96608 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96928 35308
rect 96608 33740 96928 35252
rect 96608 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96928 33740
rect 96608 32172 96928 33684
rect 96608 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96928 32172
rect 96608 30604 96928 32116
rect 96608 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96928 30604
rect 96608 29036 96928 30548
rect 96608 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96928 29036
rect 96608 27468 96928 28980
rect 96608 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96928 27468
rect 96608 25900 96928 27412
rect 96608 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96928 25900
rect 96608 24332 96928 25844
rect 96608 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96928 24332
rect 96608 22764 96928 24276
rect 96608 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96928 22764
rect 96608 21196 96928 22708
rect 96608 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96928 21196
rect 96608 19628 96928 21140
rect 96608 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96928 19628
rect 96608 18060 96928 19572
rect 96608 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96928 18060
rect 96608 16492 96928 18004
rect 96608 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96928 16492
rect 96608 14924 96928 16436
rect 96608 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96928 14924
rect 96608 13356 96928 14868
rect 111968 116060 112288 116876
rect 111968 116004 111996 116060
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 112260 116004 112288 116060
rect 111968 114492 112288 116004
rect 111968 114436 111996 114492
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 112260 114436 112288 114492
rect 111968 112924 112288 114436
rect 111968 112868 111996 112924
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 112260 112868 112288 112924
rect 111968 111356 112288 112868
rect 111968 111300 111996 111356
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 112260 111300 112288 111356
rect 111968 109788 112288 111300
rect 111968 109732 111996 109788
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 112260 109732 112288 109788
rect 111968 108220 112288 109732
rect 111968 108164 111996 108220
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 112260 108164 112288 108220
rect 111968 106652 112288 108164
rect 111968 106596 111996 106652
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 112260 106596 112288 106652
rect 111968 105084 112288 106596
rect 111968 105028 111996 105084
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 112260 105028 112288 105084
rect 111968 103516 112288 105028
rect 111968 103460 111996 103516
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 112260 103460 112288 103516
rect 111968 101948 112288 103460
rect 111968 101892 111996 101948
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 112260 101892 112288 101948
rect 111968 100380 112288 101892
rect 111968 100324 111996 100380
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 112260 100324 112288 100380
rect 111968 98812 112288 100324
rect 111968 98756 111996 98812
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 112260 98756 112288 98812
rect 111968 97244 112288 98756
rect 111968 97188 111996 97244
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 112260 97188 112288 97244
rect 111968 95676 112288 97188
rect 111968 95620 111996 95676
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 112260 95620 112288 95676
rect 111968 94108 112288 95620
rect 111968 94052 111996 94108
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 112260 94052 112288 94108
rect 111968 92540 112288 94052
rect 111968 92484 111996 92540
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 112260 92484 112288 92540
rect 111968 90972 112288 92484
rect 111968 90916 111996 90972
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 112260 90916 112288 90972
rect 111968 89404 112288 90916
rect 111968 89348 111996 89404
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 112260 89348 112288 89404
rect 111968 87836 112288 89348
rect 111968 87780 111996 87836
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 112260 87780 112288 87836
rect 111968 86268 112288 87780
rect 111968 86212 111996 86268
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 112260 86212 112288 86268
rect 111968 84700 112288 86212
rect 111968 84644 111996 84700
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 112260 84644 112288 84700
rect 111968 83132 112288 84644
rect 111968 83076 111996 83132
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 112260 83076 112288 83132
rect 111968 81564 112288 83076
rect 111968 81508 111996 81564
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 112260 81508 112288 81564
rect 111968 79996 112288 81508
rect 111968 79940 111996 79996
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 112260 79940 112288 79996
rect 111968 78428 112288 79940
rect 111968 78372 111996 78428
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 112260 78372 112288 78428
rect 111968 76860 112288 78372
rect 111968 76804 111996 76860
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 112260 76804 112288 76860
rect 111968 75292 112288 76804
rect 111968 75236 111996 75292
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 112260 75236 112288 75292
rect 111968 73724 112288 75236
rect 111968 73668 111996 73724
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 112260 73668 112288 73724
rect 111968 72156 112288 73668
rect 111968 72100 111996 72156
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 112260 72100 112288 72156
rect 111968 70588 112288 72100
rect 111968 70532 111996 70588
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 112260 70532 112288 70588
rect 111968 69020 112288 70532
rect 111968 68964 111996 69020
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 112260 68964 112288 69020
rect 111968 67452 112288 68964
rect 111968 67396 111996 67452
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 112260 67396 112288 67452
rect 111968 65884 112288 67396
rect 111968 65828 111996 65884
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 112260 65828 112288 65884
rect 111968 64316 112288 65828
rect 111968 64260 111996 64316
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 112260 64260 112288 64316
rect 111968 62748 112288 64260
rect 111968 62692 111996 62748
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 112260 62692 112288 62748
rect 111968 61180 112288 62692
rect 111968 61124 111996 61180
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 112260 61124 112288 61180
rect 111968 59612 112288 61124
rect 111968 59556 111996 59612
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 112260 59556 112288 59612
rect 111968 58044 112288 59556
rect 111968 57988 111996 58044
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 112260 57988 112288 58044
rect 111968 56476 112288 57988
rect 111968 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112288 56476
rect 111968 54908 112288 56420
rect 111968 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112288 54908
rect 111968 53340 112288 54852
rect 111968 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112288 53340
rect 111968 51772 112288 53284
rect 111968 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112288 51772
rect 111968 50204 112288 51716
rect 111968 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112288 50204
rect 111968 48636 112288 50148
rect 111968 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112288 48636
rect 111968 47068 112288 48580
rect 111968 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112288 47068
rect 111968 45500 112288 47012
rect 111968 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112288 45500
rect 111968 43932 112288 45444
rect 111968 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112288 43932
rect 111968 42364 112288 43876
rect 111968 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112288 42364
rect 111968 40796 112288 42308
rect 111968 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112288 40796
rect 111968 39228 112288 40740
rect 111968 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112288 39228
rect 111968 37660 112288 39172
rect 111968 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112288 37660
rect 111968 36092 112288 37604
rect 111968 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112288 36092
rect 111968 34524 112288 36036
rect 111968 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112288 34524
rect 111968 32956 112288 34468
rect 111968 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112288 32956
rect 111968 31388 112288 32900
rect 111968 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112288 31388
rect 111968 29820 112288 31332
rect 111968 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112288 29820
rect 111968 28252 112288 29764
rect 111968 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112288 28252
rect 111968 26684 112288 28196
rect 111968 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112288 26684
rect 111968 25116 112288 26628
rect 127328 116844 127648 116876
rect 127328 116788 127356 116844
rect 127412 116788 127460 116844
rect 127516 116788 127564 116844
rect 127620 116788 127648 116844
rect 127328 115276 127648 116788
rect 127328 115220 127356 115276
rect 127412 115220 127460 115276
rect 127516 115220 127564 115276
rect 127620 115220 127648 115276
rect 127328 113708 127648 115220
rect 127328 113652 127356 113708
rect 127412 113652 127460 113708
rect 127516 113652 127564 113708
rect 127620 113652 127648 113708
rect 127328 112140 127648 113652
rect 127328 112084 127356 112140
rect 127412 112084 127460 112140
rect 127516 112084 127564 112140
rect 127620 112084 127648 112140
rect 127328 110572 127648 112084
rect 127328 110516 127356 110572
rect 127412 110516 127460 110572
rect 127516 110516 127564 110572
rect 127620 110516 127648 110572
rect 127328 109004 127648 110516
rect 127328 108948 127356 109004
rect 127412 108948 127460 109004
rect 127516 108948 127564 109004
rect 127620 108948 127648 109004
rect 127328 107436 127648 108948
rect 127328 107380 127356 107436
rect 127412 107380 127460 107436
rect 127516 107380 127564 107436
rect 127620 107380 127648 107436
rect 127328 105868 127648 107380
rect 127328 105812 127356 105868
rect 127412 105812 127460 105868
rect 127516 105812 127564 105868
rect 127620 105812 127648 105868
rect 127328 104300 127648 105812
rect 127328 104244 127356 104300
rect 127412 104244 127460 104300
rect 127516 104244 127564 104300
rect 127620 104244 127648 104300
rect 127328 102732 127648 104244
rect 127328 102676 127356 102732
rect 127412 102676 127460 102732
rect 127516 102676 127564 102732
rect 127620 102676 127648 102732
rect 127328 101164 127648 102676
rect 127328 101108 127356 101164
rect 127412 101108 127460 101164
rect 127516 101108 127564 101164
rect 127620 101108 127648 101164
rect 127328 99596 127648 101108
rect 127328 99540 127356 99596
rect 127412 99540 127460 99596
rect 127516 99540 127564 99596
rect 127620 99540 127648 99596
rect 127328 98028 127648 99540
rect 127328 97972 127356 98028
rect 127412 97972 127460 98028
rect 127516 97972 127564 98028
rect 127620 97972 127648 98028
rect 127328 96460 127648 97972
rect 127328 96404 127356 96460
rect 127412 96404 127460 96460
rect 127516 96404 127564 96460
rect 127620 96404 127648 96460
rect 127328 94892 127648 96404
rect 127328 94836 127356 94892
rect 127412 94836 127460 94892
rect 127516 94836 127564 94892
rect 127620 94836 127648 94892
rect 127328 93324 127648 94836
rect 127328 93268 127356 93324
rect 127412 93268 127460 93324
rect 127516 93268 127564 93324
rect 127620 93268 127648 93324
rect 127328 91756 127648 93268
rect 127328 91700 127356 91756
rect 127412 91700 127460 91756
rect 127516 91700 127564 91756
rect 127620 91700 127648 91756
rect 127328 90188 127648 91700
rect 127328 90132 127356 90188
rect 127412 90132 127460 90188
rect 127516 90132 127564 90188
rect 127620 90132 127648 90188
rect 127328 88620 127648 90132
rect 127328 88564 127356 88620
rect 127412 88564 127460 88620
rect 127516 88564 127564 88620
rect 127620 88564 127648 88620
rect 127328 87052 127648 88564
rect 127328 86996 127356 87052
rect 127412 86996 127460 87052
rect 127516 86996 127564 87052
rect 127620 86996 127648 87052
rect 127328 85484 127648 86996
rect 127328 85428 127356 85484
rect 127412 85428 127460 85484
rect 127516 85428 127564 85484
rect 127620 85428 127648 85484
rect 127328 83916 127648 85428
rect 127328 83860 127356 83916
rect 127412 83860 127460 83916
rect 127516 83860 127564 83916
rect 127620 83860 127648 83916
rect 127328 82348 127648 83860
rect 127328 82292 127356 82348
rect 127412 82292 127460 82348
rect 127516 82292 127564 82348
rect 127620 82292 127648 82348
rect 127328 80780 127648 82292
rect 127328 80724 127356 80780
rect 127412 80724 127460 80780
rect 127516 80724 127564 80780
rect 127620 80724 127648 80780
rect 127328 79212 127648 80724
rect 127328 79156 127356 79212
rect 127412 79156 127460 79212
rect 127516 79156 127564 79212
rect 127620 79156 127648 79212
rect 127328 77644 127648 79156
rect 127328 77588 127356 77644
rect 127412 77588 127460 77644
rect 127516 77588 127564 77644
rect 127620 77588 127648 77644
rect 127328 76076 127648 77588
rect 127328 76020 127356 76076
rect 127412 76020 127460 76076
rect 127516 76020 127564 76076
rect 127620 76020 127648 76076
rect 127328 74508 127648 76020
rect 127328 74452 127356 74508
rect 127412 74452 127460 74508
rect 127516 74452 127564 74508
rect 127620 74452 127648 74508
rect 127328 72940 127648 74452
rect 127328 72884 127356 72940
rect 127412 72884 127460 72940
rect 127516 72884 127564 72940
rect 127620 72884 127648 72940
rect 127328 71372 127648 72884
rect 127328 71316 127356 71372
rect 127412 71316 127460 71372
rect 127516 71316 127564 71372
rect 127620 71316 127648 71372
rect 127328 69804 127648 71316
rect 127328 69748 127356 69804
rect 127412 69748 127460 69804
rect 127516 69748 127564 69804
rect 127620 69748 127648 69804
rect 127328 68236 127648 69748
rect 127328 68180 127356 68236
rect 127412 68180 127460 68236
rect 127516 68180 127564 68236
rect 127620 68180 127648 68236
rect 127328 66668 127648 68180
rect 127328 66612 127356 66668
rect 127412 66612 127460 66668
rect 127516 66612 127564 66668
rect 127620 66612 127648 66668
rect 127328 65100 127648 66612
rect 127328 65044 127356 65100
rect 127412 65044 127460 65100
rect 127516 65044 127564 65100
rect 127620 65044 127648 65100
rect 127328 63532 127648 65044
rect 127328 63476 127356 63532
rect 127412 63476 127460 63532
rect 127516 63476 127564 63532
rect 127620 63476 127648 63532
rect 127328 61964 127648 63476
rect 127328 61908 127356 61964
rect 127412 61908 127460 61964
rect 127516 61908 127564 61964
rect 127620 61908 127648 61964
rect 127328 60396 127648 61908
rect 127328 60340 127356 60396
rect 127412 60340 127460 60396
rect 127516 60340 127564 60396
rect 127620 60340 127648 60396
rect 127328 58828 127648 60340
rect 127328 58772 127356 58828
rect 127412 58772 127460 58828
rect 127516 58772 127564 58828
rect 127620 58772 127648 58828
rect 127328 57260 127648 58772
rect 127328 57204 127356 57260
rect 127412 57204 127460 57260
rect 127516 57204 127564 57260
rect 127620 57204 127648 57260
rect 127328 55692 127648 57204
rect 127328 55636 127356 55692
rect 127412 55636 127460 55692
rect 127516 55636 127564 55692
rect 127620 55636 127648 55692
rect 127328 54124 127648 55636
rect 127328 54068 127356 54124
rect 127412 54068 127460 54124
rect 127516 54068 127564 54124
rect 127620 54068 127648 54124
rect 127328 52556 127648 54068
rect 127328 52500 127356 52556
rect 127412 52500 127460 52556
rect 127516 52500 127564 52556
rect 127620 52500 127648 52556
rect 127328 50988 127648 52500
rect 127328 50932 127356 50988
rect 127412 50932 127460 50988
rect 127516 50932 127564 50988
rect 127620 50932 127648 50988
rect 127328 49420 127648 50932
rect 127328 49364 127356 49420
rect 127412 49364 127460 49420
rect 127516 49364 127564 49420
rect 127620 49364 127648 49420
rect 127328 47852 127648 49364
rect 127328 47796 127356 47852
rect 127412 47796 127460 47852
rect 127516 47796 127564 47852
rect 127620 47796 127648 47852
rect 127328 46284 127648 47796
rect 127328 46228 127356 46284
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127620 46228 127648 46284
rect 127328 44716 127648 46228
rect 127328 44660 127356 44716
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127620 44660 127648 44716
rect 127328 43148 127648 44660
rect 127328 43092 127356 43148
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127620 43092 127648 43148
rect 127328 41580 127648 43092
rect 127328 41524 127356 41580
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127620 41524 127648 41580
rect 127328 40012 127648 41524
rect 127328 39956 127356 40012
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127620 39956 127648 40012
rect 127328 38444 127648 39956
rect 127328 38388 127356 38444
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127620 38388 127648 38444
rect 127328 36876 127648 38388
rect 127328 36820 127356 36876
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127620 36820 127648 36876
rect 127328 35308 127648 36820
rect 127328 35252 127356 35308
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127620 35252 127648 35308
rect 127328 33740 127648 35252
rect 127328 33684 127356 33740
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127620 33684 127648 33740
rect 127328 32172 127648 33684
rect 127328 32116 127356 32172
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127620 32116 127648 32172
rect 127328 30604 127648 32116
rect 127328 30548 127356 30604
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127620 30548 127648 30604
rect 127328 29036 127648 30548
rect 127328 28980 127356 29036
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127620 28980 127648 29036
rect 127328 27468 127648 28980
rect 127328 27412 127356 27468
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127620 27412 127648 27468
rect 127328 25900 127648 27412
rect 127328 25844 127356 25900
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127620 25844 127648 25900
rect 111968 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112288 25116
rect 111968 23548 112288 25060
rect 111968 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112288 23548
rect 111968 21980 112288 23492
rect 124236 25396 124292 25406
rect 111968 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112288 21980
rect 111968 20412 112288 21924
rect 111968 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112288 20412
rect 111968 18844 112288 20356
rect 111968 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112288 18844
rect 111968 17276 112288 18788
rect 111968 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112288 17276
rect 111968 15708 112288 17220
rect 111968 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112288 15708
rect 111968 14140 112288 15652
rect 113148 22932 113204 22942
rect 113148 15148 113204 22876
rect 123676 20580 123732 20590
rect 121212 16996 121268 17006
rect 113148 15092 113316 15148
rect 111804 14084 111860 14094
rect 111804 13636 111860 14028
rect 111804 13570 111860 13580
rect 111968 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112288 14140
rect 96608 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96928 13356
rect 96608 11788 96928 13300
rect 96608 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96928 11788
rect 96608 10220 96928 11732
rect 111968 12572 112288 14084
rect 111968 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112288 12572
rect 96608 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96928 10220
rect 97020 11620 97076 11630
rect 97020 10276 97076 11564
rect 99820 11172 99876 11182
rect 99484 11060 99540 11070
rect 99484 10388 99540 11004
rect 99484 10322 99540 10332
rect 99708 10500 99764 10510
rect 97020 10210 97076 10220
rect 99596 10276 99652 10286
rect 99708 10276 99764 10444
rect 99652 10220 99764 10276
rect 99596 10210 99652 10220
rect 96348 10052 96404 10062
rect 95676 8484 95732 8494
rect 95676 7588 95732 8428
rect 95676 7522 95732 7532
rect 96124 7924 96180 7934
rect 96124 7364 96180 7868
rect 96124 7298 96180 7308
rect 95340 5170 95396 5180
rect 96348 5124 96404 9996
rect 96348 5058 96404 5068
rect 96608 8652 96928 10164
rect 96608 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96928 8652
rect 96608 7084 96928 8596
rect 96608 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96928 7084
rect 96608 5516 96928 7028
rect 96608 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96928 5516
rect 91420 4900 91476 4910
rect 91308 4844 91420 4900
rect 91308 4676 91364 4844
rect 91420 4834 91476 4844
rect 91308 4610 91364 4620
rect 85596 4274 85652 4284
rect 81248 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81568 3164
rect 81248 3076 81568 3108
rect 96608 3948 96928 5460
rect 99820 5236 99876 11116
rect 111968 11004 112288 12516
rect 111968 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112288 11004
rect 109788 10388 109844 10398
rect 109340 10332 109788 10388
rect 109340 10276 109396 10332
rect 109788 10322 109844 10332
rect 109340 10210 109396 10220
rect 106764 10052 106820 10062
rect 104188 9604 104244 9614
rect 99820 5170 99876 5180
rect 102172 8708 102228 8718
rect 102172 4340 102228 8652
rect 102396 8372 102452 8382
rect 102396 8036 102452 8316
rect 102396 5684 102452 7980
rect 102396 5618 102452 5628
rect 104188 6692 104244 9548
rect 104188 4452 104244 6636
rect 106764 6692 106820 9996
rect 106764 6626 106820 6636
rect 111968 9436 112288 10948
rect 111968 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112288 9436
rect 111968 7868 112288 9380
rect 111968 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112288 7868
rect 111968 6300 112288 7812
rect 111968 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112288 6300
rect 111804 5012 111860 5022
rect 111804 4788 111860 4956
rect 111804 4722 111860 4732
rect 111968 4732 112288 6244
rect 104188 4386 104244 4396
rect 111968 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112288 4732
rect 102172 4274 102228 4284
rect 96608 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96928 3948
rect 96608 3076 96928 3892
rect 111968 3164 112288 4676
rect 113260 11172 113316 15092
rect 113260 4564 113316 11116
rect 114716 11172 114772 11182
rect 114492 10164 114548 10174
rect 113932 9828 113988 9838
rect 113932 7252 113988 9772
rect 113932 4788 113988 7196
rect 113932 4722 113988 4732
rect 113260 4498 113316 4508
rect 114492 4228 114548 10108
rect 114716 7252 114772 11116
rect 114716 7186 114772 7196
rect 117292 10500 117348 10510
rect 116396 6244 116452 6254
rect 116396 5796 116452 6188
rect 116396 5730 116452 5740
rect 114492 4162 114548 4172
rect 117292 4564 117348 10444
rect 119756 9828 119812 9838
rect 119756 5124 119812 9772
rect 119756 5058 119812 5068
rect 121212 9268 121268 16940
rect 111968 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112288 3164
rect 111968 3076 112288 3108
rect 117292 2996 117348 4508
rect 121212 3556 121268 9212
rect 121324 7700 121380 7710
rect 121324 4340 121380 7644
rect 122108 6804 122164 6814
rect 122108 5012 122164 6748
rect 123676 6020 123732 20524
rect 123676 5954 123732 5964
rect 122108 4946 122164 4956
rect 121324 4274 121380 4284
rect 121772 3892 121828 3902
rect 121548 3780 121604 3790
rect 121772 3780 121828 3836
rect 121604 3724 121828 3780
rect 121548 3714 121604 3724
rect 121212 3490 121268 3500
rect 124236 3332 124292 25340
rect 124236 3266 124292 3276
rect 127328 24332 127648 25844
rect 142688 116060 143008 116876
rect 142688 116004 142716 116060
rect 142772 116004 142820 116060
rect 142876 116004 142924 116060
rect 142980 116004 143008 116060
rect 142688 114492 143008 116004
rect 142688 114436 142716 114492
rect 142772 114436 142820 114492
rect 142876 114436 142924 114492
rect 142980 114436 143008 114492
rect 142688 112924 143008 114436
rect 142688 112868 142716 112924
rect 142772 112868 142820 112924
rect 142876 112868 142924 112924
rect 142980 112868 143008 112924
rect 142688 111356 143008 112868
rect 142688 111300 142716 111356
rect 142772 111300 142820 111356
rect 142876 111300 142924 111356
rect 142980 111300 143008 111356
rect 142688 109788 143008 111300
rect 142688 109732 142716 109788
rect 142772 109732 142820 109788
rect 142876 109732 142924 109788
rect 142980 109732 143008 109788
rect 142688 108220 143008 109732
rect 142688 108164 142716 108220
rect 142772 108164 142820 108220
rect 142876 108164 142924 108220
rect 142980 108164 143008 108220
rect 142688 106652 143008 108164
rect 142688 106596 142716 106652
rect 142772 106596 142820 106652
rect 142876 106596 142924 106652
rect 142980 106596 143008 106652
rect 142688 105084 143008 106596
rect 142688 105028 142716 105084
rect 142772 105028 142820 105084
rect 142876 105028 142924 105084
rect 142980 105028 143008 105084
rect 142688 103516 143008 105028
rect 142688 103460 142716 103516
rect 142772 103460 142820 103516
rect 142876 103460 142924 103516
rect 142980 103460 143008 103516
rect 142688 101948 143008 103460
rect 142688 101892 142716 101948
rect 142772 101892 142820 101948
rect 142876 101892 142924 101948
rect 142980 101892 143008 101948
rect 142688 100380 143008 101892
rect 142688 100324 142716 100380
rect 142772 100324 142820 100380
rect 142876 100324 142924 100380
rect 142980 100324 143008 100380
rect 142688 98812 143008 100324
rect 142688 98756 142716 98812
rect 142772 98756 142820 98812
rect 142876 98756 142924 98812
rect 142980 98756 143008 98812
rect 142688 97244 143008 98756
rect 142688 97188 142716 97244
rect 142772 97188 142820 97244
rect 142876 97188 142924 97244
rect 142980 97188 143008 97244
rect 142688 95676 143008 97188
rect 142688 95620 142716 95676
rect 142772 95620 142820 95676
rect 142876 95620 142924 95676
rect 142980 95620 143008 95676
rect 142688 94108 143008 95620
rect 142688 94052 142716 94108
rect 142772 94052 142820 94108
rect 142876 94052 142924 94108
rect 142980 94052 143008 94108
rect 142688 92540 143008 94052
rect 142688 92484 142716 92540
rect 142772 92484 142820 92540
rect 142876 92484 142924 92540
rect 142980 92484 143008 92540
rect 142688 90972 143008 92484
rect 142688 90916 142716 90972
rect 142772 90916 142820 90972
rect 142876 90916 142924 90972
rect 142980 90916 143008 90972
rect 142688 89404 143008 90916
rect 142688 89348 142716 89404
rect 142772 89348 142820 89404
rect 142876 89348 142924 89404
rect 142980 89348 143008 89404
rect 142688 87836 143008 89348
rect 142688 87780 142716 87836
rect 142772 87780 142820 87836
rect 142876 87780 142924 87836
rect 142980 87780 143008 87836
rect 142688 86268 143008 87780
rect 142688 86212 142716 86268
rect 142772 86212 142820 86268
rect 142876 86212 142924 86268
rect 142980 86212 143008 86268
rect 142688 84700 143008 86212
rect 142688 84644 142716 84700
rect 142772 84644 142820 84700
rect 142876 84644 142924 84700
rect 142980 84644 143008 84700
rect 142688 83132 143008 84644
rect 142688 83076 142716 83132
rect 142772 83076 142820 83132
rect 142876 83076 142924 83132
rect 142980 83076 143008 83132
rect 142688 81564 143008 83076
rect 142688 81508 142716 81564
rect 142772 81508 142820 81564
rect 142876 81508 142924 81564
rect 142980 81508 143008 81564
rect 142688 79996 143008 81508
rect 142688 79940 142716 79996
rect 142772 79940 142820 79996
rect 142876 79940 142924 79996
rect 142980 79940 143008 79996
rect 142688 78428 143008 79940
rect 142688 78372 142716 78428
rect 142772 78372 142820 78428
rect 142876 78372 142924 78428
rect 142980 78372 143008 78428
rect 142688 76860 143008 78372
rect 142688 76804 142716 76860
rect 142772 76804 142820 76860
rect 142876 76804 142924 76860
rect 142980 76804 143008 76860
rect 142688 75292 143008 76804
rect 142688 75236 142716 75292
rect 142772 75236 142820 75292
rect 142876 75236 142924 75292
rect 142980 75236 143008 75292
rect 142688 73724 143008 75236
rect 142688 73668 142716 73724
rect 142772 73668 142820 73724
rect 142876 73668 142924 73724
rect 142980 73668 143008 73724
rect 142688 72156 143008 73668
rect 142688 72100 142716 72156
rect 142772 72100 142820 72156
rect 142876 72100 142924 72156
rect 142980 72100 143008 72156
rect 142688 70588 143008 72100
rect 142688 70532 142716 70588
rect 142772 70532 142820 70588
rect 142876 70532 142924 70588
rect 142980 70532 143008 70588
rect 142688 69020 143008 70532
rect 142688 68964 142716 69020
rect 142772 68964 142820 69020
rect 142876 68964 142924 69020
rect 142980 68964 143008 69020
rect 142688 67452 143008 68964
rect 142688 67396 142716 67452
rect 142772 67396 142820 67452
rect 142876 67396 142924 67452
rect 142980 67396 143008 67452
rect 142688 65884 143008 67396
rect 142688 65828 142716 65884
rect 142772 65828 142820 65884
rect 142876 65828 142924 65884
rect 142980 65828 143008 65884
rect 142688 64316 143008 65828
rect 142688 64260 142716 64316
rect 142772 64260 142820 64316
rect 142876 64260 142924 64316
rect 142980 64260 143008 64316
rect 142688 62748 143008 64260
rect 142688 62692 142716 62748
rect 142772 62692 142820 62748
rect 142876 62692 142924 62748
rect 142980 62692 143008 62748
rect 142688 61180 143008 62692
rect 142688 61124 142716 61180
rect 142772 61124 142820 61180
rect 142876 61124 142924 61180
rect 142980 61124 143008 61180
rect 142688 59612 143008 61124
rect 142688 59556 142716 59612
rect 142772 59556 142820 59612
rect 142876 59556 142924 59612
rect 142980 59556 143008 59612
rect 142688 58044 143008 59556
rect 142688 57988 142716 58044
rect 142772 57988 142820 58044
rect 142876 57988 142924 58044
rect 142980 57988 143008 58044
rect 142688 56476 143008 57988
rect 142688 56420 142716 56476
rect 142772 56420 142820 56476
rect 142876 56420 142924 56476
rect 142980 56420 143008 56476
rect 142688 54908 143008 56420
rect 142688 54852 142716 54908
rect 142772 54852 142820 54908
rect 142876 54852 142924 54908
rect 142980 54852 143008 54908
rect 142688 53340 143008 54852
rect 142688 53284 142716 53340
rect 142772 53284 142820 53340
rect 142876 53284 142924 53340
rect 142980 53284 143008 53340
rect 142688 51772 143008 53284
rect 142688 51716 142716 51772
rect 142772 51716 142820 51772
rect 142876 51716 142924 51772
rect 142980 51716 143008 51772
rect 142688 50204 143008 51716
rect 142688 50148 142716 50204
rect 142772 50148 142820 50204
rect 142876 50148 142924 50204
rect 142980 50148 143008 50204
rect 142688 48636 143008 50148
rect 142688 48580 142716 48636
rect 142772 48580 142820 48636
rect 142876 48580 142924 48636
rect 142980 48580 143008 48636
rect 142688 47068 143008 48580
rect 142688 47012 142716 47068
rect 142772 47012 142820 47068
rect 142876 47012 142924 47068
rect 142980 47012 143008 47068
rect 142688 45500 143008 47012
rect 142688 45444 142716 45500
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142980 45444 143008 45500
rect 142688 43932 143008 45444
rect 142688 43876 142716 43932
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142980 43876 143008 43932
rect 142688 42364 143008 43876
rect 142688 42308 142716 42364
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142980 42308 143008 42364
rect 142688 40796 143008 42308
rect 142688 40740 142716 40796
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142980 40740 143008 40796
rect 142688 39228 143008 40740
rect 142688 39172 142716 39228
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142980 39172 143008 39228
rect 142688 37660 143008 39172
rect 142688 37604 142716 37660
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142980 37604 143008 37660
rect 142688 36092 143008 37604
rect 142688 36036 142716 36092
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142980 36036 143008 36092
rect 142688 34524 143008 36036
rect 142688 34468 142716 34524
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142980 34468 143008 34524
rect 142688 32956 143008 34468
rect 142688 32900 142716 32956
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142980 32900 143008 32956
rect 142688 31388 143008 32900
rect 142688 31332 142716 31388
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142980 31332 143008 31388
rect 142688 29820 143008 31332
rect 142688 29764 142716 29820
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142980 29764 143008 29820
rect 142688 28252 143008 29764
rect 142688 28196 142716 28252
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142980 28196 143008 28252
rect 142688 26684 143008 28196
rect 142688 26628 142716 26684
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142980 26628 143008 26684
rect 127328 24276 127356 24332
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127620 24276 127648 24332
rect 127328 22764 127648 24276
rect 127328 22708 127356 22764
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127620 22708 127648 22764
rect 127328 21196 127648 22708
rect 127328 21140 127356 21196
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127620 21140 127648 21196
rect 127328 19628 127648 21140
rect 127328 19572 127356 19628
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127620 19572 127648 19628
rect 127328 18060 127648 19572
rect 127328 18004 127356 18060
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127620 18004 127648 18060
rect 127328 16492 127648 18004
rect 127328 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127648 16492
rect 127328 14924 127648 16436
rect 127328 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127648 14924
rect 127328 13356 127648 14868
rect 127328 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127648 13356
rect 127328 11788 127648 13300
rect 127328 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127648 11788
rect 127328 10220 127648 11732
rect 127328 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127648 10220
rect 127328 8652 127648 10164
rect 127328 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127648 8652
rect 127328 7084 127648 8596
rect 127328 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127648 7084
rect 127328 5516 127648 7028
rect 127328 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127648 5516
rect 127328 3948 127648 5460
rect 127708 25284 127764 25294
rect 127708 4564 127764 25228
rect 142688 25116 143008 26628
rect 142688 25060 142716 25116
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142980 25060 143008 25116
rect 142688 23548 143008 25060
rect 142688 23492 142716 23548
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142980 23492 143008 23548
rect 142688 21980 143008 23492
rect 142688 21924 142716 21980
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142980 21924 143008 21980
rect 142688 20412 143008 21924
rect 142688 20356 142716 20412
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142980 20356 143008 20412
rect 142688 18844 143008 20356
rect 142688 18788 142716 18844
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142980 18788 143008 18844
rect 142688 17276 143008 18788
rect 142688 17220 142716 17276
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142980 17220 143008 17276
rect 142688 15708 143008 17220
rect 142688 15652 142716 15708
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142980 15652 143008 15708
rect 127708 4498 127764 4508
rect 128156 15316 128212 15326
rect 127328 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127648 3948
rect 127328 3076 127648 3892
rect 128156 3332 128212 15260
rect 137004 15204 137060 15214
rect 135660 10164 135716 10174
rect 132972 6244 133028 6254
rect 132972 3780 133028 6188
rect 134652 5908 134708 5918
rect 133868 5460 133924 5470
rect 133868 4228 133924 5404
rect 133868 4162 133924 4172
rect 134652 4228 134708 5852
rect 135660 5684 135716 10108
rect 136668 8260 136724 8270
rect 136668 6580 136724 8204
rect 136668 5796 136724 6524
rect 137004 6132 137060 15148
rect 142688 14140 143008 15652
rect 142688 14084 142716 14140
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142980 14084 143008 14140
rect 142688 12572 143008 14084
rect 142688 12516 142716 12572
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142980 12516 143008 12572
rect 142688 11004 143008 12516
rect 142688 10948 142716 11004
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142980 10948 143008 11004
rect 142688 9436 143008 10948
rect 142688 9380 142716 9436
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142980 9380 143008 9436
rect 142688 7868 143008 9380
rect 142688 7812 142716 7868
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142980 7812 143008 7868
rect 140476 7364 140532 7374
rect 137340 7028 137396 7038
rect 137340 6244 137396 6972
rect 137340 6178 137396 6188
rect 137564 6804 137620 6814
rect 137004 6066 137060 6076
rect 136668 5730 136724 5740
rect 135660 4564 135716 5628
rect 135660 4498 135716 4508
rect 135884 5460 135940 5470
rect 135884 4564 135940 5404
rect 135884 4498 135940 4508
rect 134652 4162 134708 4172
rect 137564 4004 137620 6748
rect 140476 4116 140532 7308
rect 140476 4050 140532 4060
rect 142688 6300 143008 7812
rect 142688 6244 142716 6300
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142980 6244 143008 6300
rect 142688 4732 143008 6244
rect 142688 4676 142716 4732
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142980 4676 143008 4732
rect 137564 3938 137620 3948
rect 132972 3714 133028 3724
rect 128156 3266 128212 3276
rect 142688 3164 143008 4676
rect 142688 3108 142716 3164
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142980 3108 143008 3164
rect 142688 3076 143008 3108
rect 158048 116844 158368 116876
rect 158048 116788 158076 116844
rect 158132 116788 158180 116844
rect 158236 116788 158284 116844
rect 158340 116788 158368 116844
rect 158048 115276 158368 116788
rect 158048 115220 158076 115276
rect 158132 115220 158180 115276
rect 158236 115220 158284 115276
rect 158340 115220 158368 115276
rect 158048 113708 158368 115220
rect 158048 113652 158076 113708
rect 158132 113652 158180 113708
rect 158236 113652 158284 113708
rect 158340 113652 158368 113708
rect 158048 112140 158368 113652
rect 158048 112084 158076 112140
rect 158132 112084 158180 112140
rect 158236 112084 158284 112140
rect 158340 112084 158368 112140
rect 158048 110572 158368 112084
rect 158048 110516 158076 110572
rect 158132 110516 158180 110572
rect 158236 110516 158284 110572
rect 158340 110516 158368 110572
rect 158048 109004 158368 110516
rect 158048 108948 158076 109004
rect 158132 108948 158180 109004
rect 158236 108948 158284 109004
rect 158340 108948 158368 109004
rect 158048 107436 158368 108948
rect 158048 107380 158076 107436
rect 158132 107380 158180 107436
rect 158236 107380 158284 107436
rect 158340 107380 158368 107436
rect 158048 105868 158368 107380
rect 158048 105812 158076 105868
rect 158132 105812 158180 105868
rect 158236 105812 158284 105868
rect 158340 105812 158368 105868
rect 158048 104300 158368 105812
rect 158048 104244 158076 104300
rect 158132 104244 158180 104300
rect 158236 104244 158284 104300
rect 158340 104244 158368 104300
rect 158048 102732 158368 104244
rect 158048 102676 158076 102732
rect 158132 102676 158180 102732
rect 158236 102676 158284 102732
rect 158340 102676 158368 102732
rect 158048 101164 158368 102676
rect 158048 101108 158076 101164
rect 158132 101108 158180 101164
rect 158236 101108 158284 101164
rect 158340 101108 158368 101164
rect 158048 99596 158368 101108
rect 158048 99540 158076 99596
rect 158132 99540 158180 99596
rect 158236 99540 158284 99596
rect 158340 99540 158368 99596
rect 158048 98028 158368 99540
rect 158048 97972 158076 98028
rect 158132 97972 158180 98028
rect 158236 97972 158284 98028
rect 158340 97972 158368 98028
rect 158048 96460 158368 97972
rect 158048 96404 158076 96460
rect 158132 96404 158180 96460
rect 158236 96404 158284 96460
rect 158340 96404 158368 96460
rect 158048 94892 158368 96404
rect 158048 94836 158076 94892
rect 158132 94836 158180 94892
rect 158236 94836 158284 94892
rect 158340 94836 158368 94892
rect 158048 93324 158368 94836
rect 158048 93268 158076 93324
rect 158132 93268 158180 93324
rect 158236 93268 158284 93324
rect 158340 93268 158368 93324
rect 158048 91756 158368 93268
rect 158048 91700 158076 91756
rect 158132 91700 158180 91756
rect 158236 91700 158284 91756
rect 158340 91700 158368 91756
rect 158048 90188 158368 91700
rect 158048 90132 158076 90188
rect 158132 90132 158180 90188
rect 158236 90132 158284 90188
rect 158340 90132 158368 90188
rect 158048 88620 158368 90132
rect 158048 88564 158076 88620
rect 158132 88564 158180 88620
rect 158236 88564 158284 88620
rect 158340 88564 158368 88620
rect 158048 87052 158368 88564
rect 158048 86996 158076 87052
rect 158132 86996 158180 87052
rect 158236 86996 158284 87052
rect 158340 86996 158368 87052
rect 158048 85484 158368 86996
rect 158048 85428 158076 85484
rect 158132 85428 158180 85484
rect 158236 85428 158284 85484
rect 158340 85428 158368 85484
rect 158048 83916 158368 85428
rect 158048 83860 158076 83916
rect 158132 83860 158180 83916
rect 158236 83860 158284 83916
rect 158340 83860 158368 83916
rect 158048 82348 158368 83860
rect 158048 82292 158076 82348
rect 158132 82292 158180 82348
rect 158236 82292 158284 82348
rect 158340 82292 158368 82348
rect 158048 80780 158368 82292
rect 158048 80724 158076 80780
rect 158132 80724 158180 80780
rect 158236 80724 158284 80780
rect 158340 80724 158368 80780
rect 158048 79212 158368 80724
rect 158048 79156 158076 79212
rect 158132 79156 158180 79212
rect 158236 79156 158284 79212
rect 158340 79156 158368 79212
rect 158048 77644 158368 79156
rect 158048 77588 158076 77644
rect 158132 77588 158180 77644
rect 158236 77588 158284 77644
rect 158340 77588 158368 77644
rect 158048 76076 158368 77588
rect 158048 76020 158076 76076
rect 158132 76020 158180 76076
rect 158236 76020 158284 76076
rect 158340 76020 158368 76076
rect 158048 74508 158368 76020
rect 158048 74452 158076 74508
rect 158132 74452 158180 74508
rect 158236 74452 158284 74508
rect 158340 74452 158368 74508
rect 158048 72940 158368 74452
rect 158048 72884 158076 72940
rect 158132 72884 158180 72940
rect 158236 72884 158284 72940
rect 158340 72884 158368 72940
rect 158048 71372 158368 72884
rect 158048 71316 158076 71372
rect 158132 71316 158180 71372
rect 158236 71316 158284 71372
rect 158340 71316 158368 71372
rect 158048 69804 158368 71316
rect 158048 69748 158076 69804
rect 158132 69748 158180 69804
rect 158236 69748 158284 69804
rect 158340 69748 158368 69804
rect 158048 68236 158368 69748
rect 158048 68180 158076 68236
rect 158132 68180 158180 68236
rect 158236 68180 158284 68236
rect 158340 68180 158368 68236
rect 158048 66668 158368 68180
rect 158048 66612 158076 66668
rect 158132 66612 158180 66668
rect 158236 66612 158284 66668
rect 158340 66612 158368 66668
rect 158048 65100 158368 66612
rect 158048 65044 158076 65100
rect 158132 65044 158180 65100
rect 158236 65044 158284 65100
rect 158340 65044 158368 65100
rect 158048 63532 158368 65044
rect 158048 63476 158076 63532
rect 158132 63476 158180 63532
rect 158236 63476 158284 63532
rect 158340 63476 158368 63532
rect 158048 61964 158368 63476
rect 158048 61908 158076 61964
rect 158132 61908 158180 61964
rect 158236 61908 158284 61964
rect 158340 61908 158368 61964
rect 158048 60396 158368 61908
rect 158048 60340 158076 60396
rect 158132 60340 158180 60396
rect 158236 60340 158284 60396
rect 158340 60340 158368 60396
rect 158048 58828 158368 60340
rect 158048 58772 158076 58828
rect 158132 58772 158180 58828
rect 158236 58772 158284 58828
rect 158340 58772 158368 58828
rect 158048 57260 158368 58772
rect 158048 57204 158076 57260
rect 158132 57204 158180 57260
rect 158236 57204 158284 57260
rect 158340 57204 158368 57260
rect 158048 55692 158368 57204
rect 158048 55636 158076 55692
rect 158132 55636 158180 55692
rect 158236 55636 158284 55692
rect 158340 55636 158368 55692
rect 158048 54124 158368 55636
rect 158048 54068 158076 54124
rect 158132 54068 158180 54124
rect 158236 54068 158284 54124
rect 158340 54068 158368 54124
rect 158048 52556 158368 54068
rect 158048 52500 158076 52556
rect 158132 52500 158180 52556
rect 158236 52500 158284 52556
rect 158340 52500 158368 52556
rect 158048 50988 158368 52500
rect 158048 50932 158076 50988
rect 158132 50932 158180 50988
rect 158236 50932 158284 50988
rect 158340 50932 158368 50988
rect 158048 49420 158368 50932
rect 158048 49364 158076 49420
rect 158132 49364 158180 49420
rect 158236 49364 158284 49420
rect 158340 49364 158368 49420
rect 158048 47852 158368 49364
rect 158048 47796 158076 47852
rect 158132 47796 158180 47852
rect 158236 47796 158284 47852
rect 158340 47796 158368 47852
rect 158048 46284 158368 47796
rect 158048 46228 158076 46284
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158340 46228 158368 46284
rect 158048 44716 158368 46228
rect 158048 44660 158076 44716
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158340 44660 158368 44716
rect 158048 43148 158368 44660
rect 158048 43092 158076 43148
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158340 43092 158368 43148
rect 158048 41580 158368 43092
rect 158048 41524 158076 41580
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158340 41524 158368 41580
rect 158048 40012 158368 41524
rect 158048 39956 158076 40012
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158340 39956 158368 40012
rect 158048 38444 158368 39956
rect 158048 38388 158076 38444
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158340 38388 158368 38444
rect 158048 36876 158368 38388
rect 158048 36820 158076 36876
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158340 36820 158368 36876
rect 158048 35308 158368 36820
rect 158048 35252 158076 35308
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158340 35252 158368 35308
rect 158048 33740 158368 35252
rect 158048 33684 158076 33740
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158340 33684 158368 33740
rect 158048 32172 158368 33684
rect 158048 32116 158076 32172
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158340 32116 158368 32172
rect 158048 30604 158368 32116
rect 158048 30548 158076 30604
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158340 30548 158368 30604
rect 158048 29036 158368 30548
rect 158048 28980 158076 29036
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158340 28980 158368 29036
rect 158048 27468 158368 28980
rect 158048 27412 158076 27468
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158340 27412 158368 27468
rect 158048 25900 158368 27412
rect 158048 25844 158076 25900
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158340 25844 158368 25900
rect 158048 24332 158368 25844
rect 158048 24276 158076 24332
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158340 24276 158368 24332
rect 158048 22764 158368 24276
rect 158048 22708 158076 22764
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158340 22708 158368 22764
rect 158048 21196 158368 22708
rect 158048 21140 158076 21196
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158340 21140 158368 21196
rect 158048 19628 158368 21140
rect 158048 19572 158076 19628
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158340 19572 158368 19628
rect 158048 18060 158368 19572
rect 158048 18004 158076 18060
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158340 18004 158368 18060
rect 158048 16492 158368 18004
rect 158048 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158368 16492
rect 158048 14924 158368 16436
rect 158048 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158368 14924
rect 158048 13356 158368 14868
rect 158048 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158368 13356
rect 158048 11788 158368 13300
rect 158048 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158368 11788
rect 158048 10220 158368 11732
rect 158048 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158368 10220
rect 158048 8652 158368 10164
rect 158048 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158368 8652
rect 158048 7084 158368 8596
rect 158048 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158368 7084
rect 158048 5516 158368 7028
rect 158048 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158368 5516
rect 158048 3948 158368 5460
rect 158048 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158368 3948
rect 158048 3076 158368 3892
rect 173408 116060 173728 116876
rect 173408 116004 173436 116060
rect 173492 116004 173540 116060
rect 173596 116004 173644 116060
rect 173700 116004 173728 116060
rect 173408 114492 173728 116004
rect 173408 114436 173436 114492
rect 173492 114436 173540 114492
rect 173596 114436 173644 114492
rect 173700 114436 173728 114492
rect 173408 112924 173728 114436
rect 173408 112868 173436 112924
rect 173492 112868 173540 112924
rect 173596 112868 173644 112924
rect 173700 112868 173728 112924
rect 173408 111356 173728 112868
rect 173408 111300 173436 111356
rect 173492 111300 173540 111356
rect 173596 111300 173644 111356
rect 173700 111300 173728 111356
rect 173408 109788 173728 111300
rect 173408 109732 173436 109788
rect 173492 109732 173540 109788
rect 173596 109732 173644 109788
rect 173700 109732 173728 109788
rect 173408 108220 173728 109732
rect 173408 108164 173436 108220
rect 173492 108164 173540 108220
rect 173596 108164 173644 108220
rect 173700 108164 173728 108220
rect 173408 106652 173728 108164
rect 173408 106596 173436 106652
rect 173492 106596 173540 106652
rect 173596 106596 173644 106652
rect 173700 106596 173728 106652
rect 173408 105084 173728 106596
rect 173408 105028 173436 105084
rect 173492 105028 173540 105084
rect 173596 105028 173644 105084
rect 173700 105028 173728 105084
rect 173408 103516 173728 105028
rect 173408 103460 173436 103516
rect 173492 103460 173540 103516
rect 173596 103460 173644 103516
rect 173700 103460 173728 103516
rect 173408 101948 173728 103460
rect 173408 101892 173436 101948
rect 173492 101892 173540 101948
rect 173596 101892 173644 101948
rect 173700 101892 173728 101948
rect 173408 100380 173728 101892
rect 173408 100324 173436 100380
rect 173492 100324 173540 100380
rect 173596 100324 173644 100380
rect 173700 100324 173728 100380
rect 173408 98812 173728 100324
rect 173408 98756 173436 98812
rect 173492 98756 173540 98812
rect 173596 98756 173644 98812
rect 173700 98756 173728 98812
rect 173408 97244 173728 98756
rect 173408 97188 173436 97244
rect 173492 97188 173540 97244
rect 173596 97188 173644 97244
rect 173700 97188 173728 97244
rect 173408 95676 173728 97188
rect 173408 95620 173436 95676
rect 173492 95620 173540 95676
rect 173596 95620 173644 95676
rect 173700 95620 173728 95676
rect 173408 94108 173728 95620
rect 173408 94052 173436 94108
rect 173492 94052 173540 94108
rect 173596 94052 173644 94108
rect 173700 94052 173728 94108
rect 173408 92540 173728 94052
rect 173408 92484 173436 92540
rect 173492 92484 173540 92540
rect 173596 92484 173644 92540
rect 173700 92484 173728 92540
rect 173408 90972 173728 92484
rect 173408 90916 173436 90972
rect 173492 90916 173540 90972
rect 173596 90916 173644 90972
rect 173700 90916 173728 90972
rect 173408 89404 173728 90916
rect 173408 89348 173436 89404
rect 173492 89348 173540 89404
rect 173596 89348 173644 89404
rect 173700 89348 173728 89404
rect 173408 87836 173728 89348
rect 173408 87780 173436 87836
rect 173492 87780 173540 87836
rect 173596 87780 173644 87836
rect 173700 87780 173728 87836
rect 173408 86268 173728 87780
rect 173408 86212 173436 86268
rect 173492 86212 173540 86268
rect 173596 86212 173644 86268
rect 173700 86212 173728 86268
rect 173408 84700 173728 86212
rect 173408 84644 173436 84700
rect 173492 84644 173540 84700
rect 173596 84644 173644 84700
rect 173700 84644 173728 84700
rect 173408 83132 173728 84644
rect 173408 83076 173436 83132
rect 173492 83076 173540 83132
rect 173596 83076 173644 83132
rect 173700 83076 173728 83132
rect 173408 81564 173728 83076
rect 173408 81508 173436 81564
rect 173492 81508 173540 81564
rect 173596 81508 173644 81564
rect 173700 81508 173728 81564
rect 173408 79996 173728 81508
rect 173408 79940 173436 79996
rect 173492 79940 173540 79996
rect 173596 79940 173644 79996
rect 173700 79940 173728 79996
rect 173408 78428 173728 79940
rect 173408 78372 173436 78428
rect 173492 78372 173540 78428
rect 173596 78372 173644 78428
rect 173700 78372 173728 78428
rect 173408 76860 173728 78372
rect 173408 76804 173436 76860
rect 173492 76804 173540 76860
rect 173596 76804 173644 76860
rect 173700 76804 173728 76860
rect 173408 75292 173728 76804
rect 173408 75236 173436 75292
rect 173492 75236 173540 75292
rect 173596 75236 173644 75292
rect 173700 75236 173728 75292
rect 173408 73724 173728 75236
rect 173408 73668 173436 73724
rect 173492 73668 173540 73724
rect 173596 73668 173644 73724
rect 173700 73668 173728 73724
rect 173408 72156 173728 73668
rect 173408 72100 173436 72156
rect 173492 72100 173540 72156
rect 173596 72100 173644 72156
rect 173700 72100 173728 72156
rect 173408 70588 173728 72100
rect 173408 70532 173436 70588
rect 173492 70532 173540 70588
rect 173596 70532 173644 70588
rect 173700 70532 173728 70588
rect 173408 69020 173728 70532
rect 173408 68964 173436 69020
rect 173492 68964 173540 69020
rect 173596 68964 173644 69020
rect 173700 68964 173728 69020
rect 173408 67452 173728 68964
rect 173408 67396 173436 67452
rect 173492 67396 173540 67452
rect 173596 67396 173644 67452
rect 173700 67396 173728 67452
rect 173408 65884 173728 67396
rect 173408 65828 173436 65884
rect 173492 65828 173540 65884
rect 173596 65828 173644 65884
rect 173700 65828 173728 65884
rect 173408 64316 173728 65828
rect 173408 64260 173436 64316
rect 173492 64260 173540 64316
rect 173596 64260 173644 64316
rect 173700 64260 173728 64316
rect 173408 62748 173728 64260
rect 173408 62692 173436 62748
rect 173492 62692 173540 62748
rect 173596 62692 173644 62748
rect 173700 62692 173728 62748
rect 173408 61180 173728 62692
rect 173408 61124 173436 61180
rect 173492 61124 173540 61180
rect 173596 61124 173644 61180
rect 173700 61124 173728 61180
rect 173408 59612 173728 61124
rect 173408 59556 173436 59612
rect 173492 59556 173540 59612
rect 173596 59556 173644 59612
rect 173700 59556 173728 59612
rect 173408 58044 173728 59556
rect 173408 57988 173436 58044
rect 173492 57988 173540 58044
rect 173596 57988 173644 58044
rect 173700 57988 173728 58044
rect 173408 56476 173728 57988
rect 173408 56420 173436 56476
rect 173492 56420 173540 56476
rect 173596 56420 173644 56476
rect 173700 56420 173728 56476
rect 173408 54908 173728 56420
rect 173408 54852 173436 54908
rect 173492 54852 173540 54908
rect 173596 54852 173644 54908
rect 173700 54852 173728 54908
rect 173408 53340 173728 54852
rect 173408 53284 173436 53340
rect 173492 53284 173540 53340
rect 173596 53284 173644 53340
rect 173700 53284 173728 53340
rect 173408 51772 173728 53284
rect 173408 51716 173436 51772
rect 173492 51716 173540 51772
rect 173596 51716 173644 51772
rect 173700 51716 173728 51772
rect 173408 50204 173728 51716
rect 173408 50148 173436 50204
rect 173492 50148 173540 50204
rect 173596 50148 173644 50204
rect 173700 50148 173728 50204
rect 173408 48636 173728 50148
rect 173408 48580 173436 48636
rect 173492 48580 173540 48636
rect 173596 48580 173644 48636
rect 173700 48580 173728 48636
rect 173408 47068 173728 48580
rect 173408 47012 173436 47068
rect 173492 47012 173540 47068
rect 173596 47012 173644 47068
rect 173700 47012 173728 47068
rect 173408 45500 173728 47012
rect 173408 45444 173436 45500
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173700 45444 173728 45500
rect 173408 43932 173728 45444
rect 173408 43876 173436 43932
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173700 43876 173728 43932
rect 173408 42364 173728 43876
rect 173408 42308 173436 42364
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173700 42308 173728 42364
rect 173408 40796 173728 42308
rect 173408 40740 173436 40796
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173700 40740 173728 40796
rect 173408 39228 173728 40740
rect 173408 39172 173436 39228
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173700 39172 173728 39228
rect 173408 37660 173728 39172
rect 173408 37604 173436 37660
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173700 37604 173728 37660
rect 173408 36092 173728 37604
rect 173408 36036 173436 36092
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173700 36036 173728 36092
rect 173408 34524 173728 36036
rect 173408 34468 173436 34524
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173700 34468 173728 34524
rect 173408 32956 173728 34468
rect 173408 32900 173436 32956
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173700 32900 173728 32956
rect 173408 31388 173728 32900
rect 173408 31332 173436 31388
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173700 31332 173728 31388
rect 173408 29820 173728 31332
rect 173408 29764 173436 29820
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173700 29764 173728 29820
rect 173408 28252 173728 29764
rect 173408 28196 173436 28252
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173700 28196 173728 28252
rect 173408 26684 173728 28196
rect 173408 26628 173436 26684
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173700 26628 173728 26684
rect 173408 25116 173728 26628
rect 173408 25060 173436 25116
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173700 25060 173728 25116
rect 173408 23548 173728 25060
rect 173408 23492 173436 23548
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173700 23492 173728 23548
rect 173408 21980 173728 23492
rect 173408 21924 173436 21980
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173700 21924 173728 21980
rect 173408 20412 173728 21924
rect 173408 20356 173436 20412
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173700 20356 173728 20412
rect 173408 18844 173728 20356
rect 173408 18788 173436 18844
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173700 18788 173728 18844
rect 173408 17276 173728 18788
rect 173408 17220 173436 17276
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173700 17220 173728 17276
rect 173408 15708 173728 17220
rect 173408 15652 173436 15708
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173700 15652 173728 15708
rect 173408 14140 173728 15652
rect 173408 14084 173436 14140
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173700 14084 173728 14140
rect 173408 12572 173728 14084
rect 173408 12516 173436 12572
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173700 12516 173728 12572
rect 173408 11004 173728 12516
rect 173408 10948 173436 11004
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173700 10948 173728 11004
rect 173408 9436 173728 10948
rect 173408 9380 173436 9436
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173700 9380 173728 9436
rect 173408 7868 173728 9380
rect 173408 7812 173436 7868
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173700 7812 173728 7868
rect 173408 6300 173728 7812
rect 173408 6244 173436 6300
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173700 6244 173728 6300
rect 173408 4732 173728 6244
rect 173408 4676 173436 4732
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173700 4676 173728 4732
rect 173408 3164 173728 4676
rect 173408 3108 173436 3164
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173700 3108 173728 3164
rect 173408 3076 173728 3108
rect 117292 2930 117348 2940
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__I pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 92064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I
timestamp 1666464484
transform 1 0 137760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I
timestamp 1666464484
transform 1 0 133840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__A2
timestamp 1666464484
transform 1 0 93072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__A1
timestamp 1666464484
transform 1 0 63728 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__A2
timestamp 1666464484
transform -1 0 61824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__I
timestamp 1666464484
transform -1 0 56112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I
timestamp 1666464484
transform -1 0 40992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__I
timestamp 1666464484
transform -1 0 35392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__I
timestamp 1666464484
transform 1 0 103600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__I
timestamp 1666464484
transform 1 0 116928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__A2
timestamp 1666464484
transform -1 0 122640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__I
timestamp 1666464484
transform 1 0 128912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A1
timestamp 1666464484
transform -1 0 130032 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A1
timestamp 1666464484
transform 1 0 124880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A2
timestamp 1666464484
transform 1 0 125328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A1
timestamp 1666464484
transform 1 0 126784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A2
timestamp 1666464484
transform 1 0 124992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__I
timestamp 1666464484
transform -1 0 141008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__A2
timestamp 1666464484
transform 1 0 96320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A2
timestamp 1666464484
transform 1 0 124208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__A1
timestamp 1666464484
transform 1 0 117824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__A2
timestamp 1666464484
transform 1 0 115024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__A3
timestamp 1666464484
transform -1 0 114576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__A1
timestamp 1666464484
transform -1 0 140112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__A2
timestamp 1666464484
transform 1 0 139888 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A1
timestamp 1666464484
transform 1 0 136080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__A1
timestamp 1666464484
transform -1 0 128688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__A1
timestamp 1666464484
transform -1 0 131152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A1
timestamp 1666464484
transform -1 0 132048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A2
timestamp 1666464484
transform -1 0 132496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__A1
timestamp 1666464484
transform 1 0 128016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__A2
timestamp 1666464484
transform 1 0 128912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__A3
timestamp 1666464484
transform -1 0 129584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A1
timestamp 1666464484
transform 1 0 127232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A2
timestamp 1666464484
transform 1 0 126448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A3
timestamp 1666464484
transform 1 0 126896 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__A2
timestamp 1666464484
transform 1 0 141680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__A2
timestamp 1666464484
transform 1 0 137200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__A2
timestamp 1666464484
transform -1 0 142352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__A2
timestamp 1666464484
transform -1 0 141008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A1
timestamp 1666464484
transform -1 0 138768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A2
timestamp 1666464484
transform 1 0 136864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A3
timestamp 1666464484
transform 1 0 137760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A4
timestamp 1666464484
transform -1 0 139216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__A2
timestamp 1666464484
transform 1 0 147728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__A2
timestamp 1666464484
transform 1 0 148736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A1
timestamp 1666464484
transform -1 0 149744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A2
timestamp 1666464484
transform 1 0 149072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__A2
timestamp 1666464484
transform -1 0 135184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A1
timestamp 1666464484
transform 1 0 139104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A2
timestamp 1666464484
transform -1 0 140560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A3
timestamp 1666464484
transform 1 0 141232 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A4
timestamp 1666464484
transform 1 0 138208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A2
timestamp 1666464484
transform 1 0 148176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__A2
timestamp 1666464484
transform -1 0 130704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A2
timestamp 1666464484
transform 1 0 146608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A1
timestamp 1666464484
transform -1 0 134176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A2
timestamp 1666464484
transform 1 0 132720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A3
timestamp 1666464484
transform 1 0 136192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A4
timestamp 1666464484
transform 1 0 134400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__A1
timestamp 1666464484
transform 1 0 143472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__A2
timestamp 1666464484
transform 1 0 146048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__B
timestamp 1666464484
transform 1 0 143920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A2
timestamp 1666464484
transform 1 0 144480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A2
timestamp 1666464484
transform 1 0 147280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__B
timestamp 1666464484
transform 1 0 145712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__A2
timestamp 1666464484
transform 1 0 138096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__A2
timestamp 1666464484
transform -1 0 142800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A2
timestamp 1666464484
transform -1 0 123872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A4
timestamp 1666464484
transform -1 0 124768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__I
timestamp 1666464484
transform 1 0 93968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A1
timestamp 1666464484
transform -1 0 32592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A2
timestamp 1666464484
transform -1 0 39648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A1
timestamp 1666464484
transform 1 0 76160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A2
timestamp 1666464484
transform 1 0 73360 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A1
timestamp 1666464484
transform -1 0 76720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__I
timestamp 1666464484
transform 1 0 57120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A1
timestamp 1666464484
transform -1 0 65632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A2
timestamp 1666464484
transform -1 0 68320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__B1
timestamp 1666464484
transform 1 0 64288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__B2
timestamp 1666464484
transform -1 0 64848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__I
timestamp 1666464484
transform 1 0 33488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__I
timestamp 1666464484
transform 1 0 36960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__A3
timestamp 1666464484
transform 1 0 32816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__A4
timestamp 1666464484
transform -1 0 41552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A1
timestamp 1666464484
transform -1 0 60032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__B
timestamp 1666464484
transform -1 0 58912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__I
timestamp 1666464484
transform 1 0 73584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__I
timestamp 1666464484
transform -1 0 74256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__I
timestamp 1666464484
transform 1 0 58352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__I
timestamp 1666464484
transform -1 0 79184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__A3
timestamp 1666464484
transform -1 0 42672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__A4
timestamp 1666464484
transform -1 0 36960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A1
timestamp 1666464484
transform -1 0 69216 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A2
timestamp 1666464484
transform -1 0 58688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__B1
timestamp 1666464484
transform -1 0 69664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__C
timestamp 1666464484
transform -1 0 60816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__A1
timestamp 1666464484
transform -1 0 67536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__A1
timestamp 1666464484
transform 1 0 66864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__I
timestamp 1666464484
transform -1 0 79744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__B
timestamp 1666464484
transform 1 0 66080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__A1
timestamp 1666464484
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__B
timestamp 1666464484
transform -1 0 77840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__A3
timestamp 1666464484
transform -1 0 42224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__A4
timestamp 1666464484
transform 1 0 42560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__A1
timestamp 1666464484
transform -1 0 70336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__A2
timestamp 1666464484
transform -1 0 71344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__B2
timestamp 1666464484
transform -1 0 70896 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__C
timestamp 1666464484
transform -1 0 61488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__A1
timestamp 1666464484
transform 1 0 66192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A1
timestamp 1666464484
transform -1 0 57344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A3
timestamp 1666464484
transform -1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A4
timestamp 1666464484
transform 1 0 43008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__A1
timestamp 1666464484
transform -1 0 70224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__A2
timestamp 1666464484
transform -1 0 69776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__B1
timestamp 1666464484
transform -1 0 61824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__C
timestamp 1666464484
transform -1 0 64064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__A1
timestamp 1666464484
transform -1 0 65520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__I
timestamp 1666464484
transform -1 0 131600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__A1
timestamp 1666464484
transform -1 0 128464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__I
timestamp 1666464484
transform 1 0 24752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A1
timestamp 1666464484
transform 1 0 67312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A2
timestamp 1666464484
transform 1 0 62944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A3
timestamp 1666464484
transform 1 0 58800 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A4
timestamp 1666464484
transform 1 0 65632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__A1
timestamp 1666464484
transform 1 0 61712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__A2
timestamp 1666464484
transform -1 0 68768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__I
timestamp 1666464484
transform -1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__A2
timestamp 1666464484
transform -1 0 64848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A1
timestamp 1666464484
transform -1 0 61936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A2
timestamp 1666464484
transform -1 0 72352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__B1
timestamp 1666464484
transform -1 0 72800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__C2
timestamp 1666464484
transform -1 0 71120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__A1
timestamp 1666464484
transform -1 0 72016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__I
timestamp 1666464484
transform 1 0 77168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A1
timestamp 1666464484
transform 1 0 70112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A2
timestamp 1666464484
transform 1 0 69664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A1
timestamp 1666464484
transform 1 0 71008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A1
timestamp 1666464484
transform -1 0 75264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A2
timestamp 1666464484
transform -1 0 74816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__C2
timestamp 1666464484
transform -1 0 73248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A1
timestamp 1666464484
transform 1 0 70000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A2
timestamp 1666464484
transform -1 0 70672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__A3
timestamp 1666464484
transform 1 0 68096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A1
timestamp 1666464484
transform 1 0 73472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__A1
timestamp 1666464484
transform -1 0 63728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__A2
timestamp 1666464484
transform -1 0 75040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__C2
timestamp 1666464484
transform -1 0 72800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__I
timestamp 1666464484
transform -1 0 135296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A2
timestamp 1666464484
transform 1 0 134288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__I
timestamp 1666464484
transform 1 0 78400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A1
timestamp 1666464484
transform 1 0 75376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A2
timestamp 1666464484
transform 1 0 70560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A3
timestamp 1666464484
transform 1 0 64624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A4
timestamp 1666464484
transform -1 0 71792 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__A1
timestamp 1666464484
transform 1 0 68544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A1
timestamp 1666464484
transform -1 0 79184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A2
timestamp 1666464484
transform -1 0 68992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__C2
timestamp 1666464484
transform -1 0 77168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__A1
timestamp 1666464484
transform -1 0 80976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__A2
timestamp 1666464484
transform 1 0 79968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A1
timestamp 1666464484
transform 1 0 82544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__I
timestamp 1666464484
transform -1 0 85568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A1
timestamp 1666464484
transform -1 0 78064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__467__A1
timestamp 1666464484
transform 1 0 80080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__A2
timestamp 1666464484
transform -1 0 80752 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A1
timestamp 1666464484
transform -1 0 83216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A2
timestamp 1666464484
transform -1 0 84896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__C2
timestamp 1666464484
transform -1 0 82320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__A2
timestamp 1666464484
transform 1 0 79184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__A1
timestamp 1666464484
transform 1 0 79632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__B
timestamp 1666464484
transform 1 0 80528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A1
timestamp 1666464484
transform 1 0 76048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A2
timestamp 1666464484
transform 1 0 76496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__A1
timestamp 1666464484
transform -1 0 77168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__A1
timestamp 1666464484
transform -1 0 86576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__A2
timestamp 1666464484
transform -1 0 87136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__B2
timestamp 1666464484
transform -1 0 84672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__I
timestamp 1666464484
transform -1 0 103376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__479__B
timestamp 1666464484
transform 1 0 86912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__I
timestamp 1666464484
transform 1 0 80976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A1
timestamp 1666464484
transform 1 0 81536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__A1
timestamp 1666464484
transform -1 0 78064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__A2
timestamp 1666464484
transform -1 0 86016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__C2
timestamp 1666464484
transform 1 0 75600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__I
timestamp 1666464484
transform 1 0 51968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__A1
timestamp 1666464484
transform -1 0 76272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__486__A1
timestamp 1666464484
transform 1 0 83664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__486__A2
timestamp 1666464484
transform 1 0 87696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__A1
timestamp 1666464484
transform -1 0 87696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__A2
timestamp 1666464484
transform -1 0 87024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__C2
timestamp 1666464484
transform -1 0 79968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A1
timestamp 1666464484
transform 1 0 86240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A2
timestamp 1666464484
transform 1 0 86688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__A1
timestamp 1666464484
transform 1 0 90832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__A1
timestamp 1666464484
transform -1 0 91616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__A2
timestamp 1666464484
transform -1 0 92064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__B1
timestamp 1666464484
transform 1 0 89152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__C2
timestamp 1666464484
transform -1 0 89376 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__A1
timestamp 1666464484
transform 1 0 89376 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A1
timestamp 1666464484
transform -1 0 89824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A1
timestamp 1666464484
transform -1 0 91840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A2
timestamp 1666464484
transform 1 0 93744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__B1
timestamp 1666464484
transform -1 0 88816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__C2
timestamp 1666464484
transform -1 0 88368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__I
timestamp 1666464484
transform 1 0 81424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__I
timestamp 1666464484
transform -1 0 67872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A1
timestamp 1666464484
transform 1 0 87696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A2
timestamp 1666464484
transform 1 0 87248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A3
timestamp 1666464484
transform 1 0 85792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A4
timestamp 1666464484
transform -1 0 80752 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__A1
timestamp 1666464484
transform 1 0 80080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A1
timestamp 1666464484
transform 1 0 81648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__B2
timestamp 1666464484
transform -1 0 81424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A3
timestamp 1666464484
transform 1 0 143024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A1
timestamp 1666464484
transform -1 0 82768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__B1
timestamp 1666464484
transform -1 0 84224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__C
timestamp 1666464484
transform -1 0 76608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A1
timestamp 1666464484
transform 1 0 82768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__I
timestamp 1666464484
transform 1 0 77168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A1
timestamp 1666464484
transform 1 0 82656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A2
timestamp 1666464484
transform 1 0 88368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A1
timestamp 1666464484
transform -1 0 93744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A2
timestamp 1666464484
transform 1 0 92288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__B1
timestamp 1666464484
transform 1 0 90048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__C2
timestamp 1666464484
transform 1 0 88144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__A1
timestamp 1666464484
transform 1 0 90384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A1
timestamp 1666464484
transform -1 0 136192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A2
timestamp 1666464484
transform -1 0 135744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__A2
timestamp 1666464484
transform -1 0 16464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__A1
timestamp 1666464484
transform -1 0 78176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__A2
timestamp 1666464484
transform 1 0 78512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A1
timestamp 1666464484
transform 1 0 74928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__I
timestamp 1666464484
transform 1 0 116704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__A1
timestamp 1666464484
transform 1 0 90944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__A2
timestamp 1666464484
transform 1 0 93072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A1
timestamp 1666464484
transform 1 0 112112 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A2
timestamp 1666464484
transform -1 0 107072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__A2
timestamp 1666464484
transform -1 0 78288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__I
timestamp 1666464484
transform -1 0 115136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A1
timestamp 1666464484
transform -1 0 123536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A2
timestamp 1666464484
transform -1 0 122528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__B2
timestamp 1666464484
transform -1 0 117824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__C2
timestamp 1666464484
transform -1 0 117376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A1
timestamp 1666464484
transform 1 0 103488 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A2
timestamp 1666464484
transform 1 0 104608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__I
timestamp 1666464484
transform 1 0 121968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A1
timestamp 1666464484
transform 1 0 107296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A2
timestamp 1666464484
transform 1 0 112560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__B
timestamp 1666464484
transform 1 0 113456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__A1
timestamp 1666464484
transform 1 0 79632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__A2
timestamp 1666464484
transform 1 0 80080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__A1
timestamp 1666464484
transform -1 0 83776 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__A2
timestamp 1666464484
transform -1 0 83328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__I
timestamp 1666464484
transform 1 0 120960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__A2
timestamp 1666464484
transform 1 0 121072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A1
timestamp 1666464484
transform -1 0 121632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A2
timestamp 1666464484
transform 1 0 127120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__B2
timestamp 1666464484
transform 1 0 120960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A1
timestamp 1666464484
transform -1 0 105280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A2
timestamp 1666464484
transform -1 0 106176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__I
timestamp 1666464484
transform -1 0 116144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__I
timestamp 1666464484
transform 1 0 113456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__A1
timestamp 1666464484
transform 1 0 121408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__I
timestamp 1666464484
transform 1 0 115360 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__A1
timestamp 1666464484
transform -1 0 125664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__A2
timestamp 1666464484
transform -1 0 123088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__C2
timestamp 1666464484
transform 1 0 121968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A1
timestamp 1666464484
transform 1 0 120064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A2
timestamp 1666464484
transform 1 0 120624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A1
timestamp 1666464484
transform 1 0 119616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__B
timestamp 1666464484
transform 1 0 119168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__A1
timestamp 1666464484
transform -1 0 123984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__A2
timestamp 1666464484
transform -1 0 122976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__B2
timestamp 1666464484
transform 1 0 119840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__A1
timestamp 1666464484
transform 1 0 122864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__A1
timestamp 1666464484
transform -1 0 126112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__A2
timestamp 1666464484
transform -1 0 123536 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__C2
timestamp 1666464484
transform 1 0 123200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__A1
timestamp 1666464484
transform 1 0 122416 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__A1
timestamp 1666464484
transform 1 0 108528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__A2
timestamp 1666464484
transform 1 0 105952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A1
timestamp 1666464484
transform 1 0 113904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A2
timestamp 1666464484
transform 1 0 114352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A3
timestamp 1666464484
transform 1 0 108976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__A1
timestamp 1666464484
transform 1 0 115472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__B
timestamp 1666464484
transform 1 0 117824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__A1
timestamp 1666464484
transform -1 0 126560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__A2
timestamp 1666464484
transform -1 0 124320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__B2
timestamp 1666464484
transform 1 0 121856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__A2
timestamp 1666464484
transform -1 0 118944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__B
timestamp 1666464484
transform 1 0 118272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__550__I
timestamp 1666464484
transform 1 0 114128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__A1
timestamp 1666464484
transform -1 0 113680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__A2
timestamp 1666464484
transform -1 0 114800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__A1
timestamp 1666464484
transform -1 0 118272 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__A2
timestamp 1666464484
transform -1 0 122080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__B1
timestamp 1666464484
transform -1 0 115360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__C2
timestamp 1666464484
transform 1 0 121520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__554__I
timestamp 1666464484
transform 1 0 108528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__A1
timestamp 1666464484
transform 1 0 143920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__A2
timestamp 1666464484
transform 1 0 142576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__A1
timestamp 1666464484
transform 1 0 113680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__A2
timestamp 1666464484
transform 1 0 117376 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__A1
timestamp 1666464484
transform 1 0 113904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__A2
timestamp 1666464484
transform 1 0 116368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__A1
timestamp 1666464484
transform -1 0 116032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__A2
timestamp 1666464484
transform -1 0 114800 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__B1
timestamp 1666464484
transform 1 0 122752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__C2
timestamp 1666464484
transform 1 0 113120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__559__A1
timestamp 1666464484
transform 1 0 116928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__A1
timestamp 1666464484
transform -1 0 17472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__A1
timestamp 1666464484
transform 1 0 79632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__A2
timestamp 1666464484
transform 1 0 79184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__A1
timestamp 1666464484
transform 1 0 80528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__563__I
timestamp 1666464484
transform 1 0 105056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__A1
timestamp 1666464484
transform 1 0 113904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__A2
timestamp 1666464484
transform -1 0 108304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__565__A1
timestamp 1666464484
transform 1 0 113680 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__A2
timestamp 1666464484
transform -1 0 79856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__I
timestamp 1666464484
transform -1 0 94528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__A1
timestamp 1666464484
transform -1 0 117152 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__A2
timestamp 1666464484
transform -1 0 114128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__B1
timestamp 1666464484
transform 1 0 113008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__C1
timestamp 1666464484
transform 1 0 116480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__C2
timestamp 1666464484
transform 1 0 113232 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__569__A1
timestamp 1666464484
transform 1 0 114800 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__570__A1
timestamp 1666464484
transform -1 0 130480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__571__I
timestamp 1666464484
transform 1 0 107520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__I
timestamp 1666464484
transform -1 0 110432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__A1
timestamp 1666464484
transform 1 0 115920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__A2
timestamp 1666464484
transform 1 0 107408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__A3
timestamp 1666464484
transform -1 0 115024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__574__I
timestamp 1666464484
transform 1 0 93744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__I
timestamp 1666464484
transform 1 0 106176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__576__A1
timestamp 1666464484
transform 1 0 104048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__576__A2
timestamp 1666464484
transform 1 0 106848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__577__A1
timestamp 1666464484
transform 1 0 111664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__577__A2
timestamp 1666464484
transform 1 0 110768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__577__A3
timestamp 1666464484
transform 1 0 110320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__I
timestamp 1666464484
transform 1 0 106400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__579__A1
timestamp 1666464484
transform 1 0 101920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A1
timestamp 1666464484
transform -1 0 107296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A2
timestamp 1666464484
transform -1 0 107520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__B2
timestamp 1666464484
transform 1 0 102368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__A1
timestamp 1666464484
transform 1 0 105728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__I
timestamp 1666464484
transform 1 0 105504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__583__A1
timestamp 1666464484
transform 1 0 105952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A1
timestamp 1666464484
transform -1 0 107184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A2
timestamp 1666464484
transform 1 0 113008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__B1
timestamp 1666464484
transform -1 0 107072 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__C1
timestamp 1666464484
transform -1 0 107520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__C2
timestamp 1666464484
transform 1 0 106400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A1
timestamp 1666464484
transform 1 0 106624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__586__I
timestamp 1666464484
transform 1 0 97216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__A1
timestamp 1666464484
transform 1 0 101472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__A2
timestamp 1666464484
transform 1 0 99904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__A3
timestamp 1666464484
transform 1 0 101024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__A1
timestamp 1666464484
transform 1 0 99008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__B
timestamp 1666464484
transform 1 0 99456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__A1
timestamp 1666464484
transform -1 0 139664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__A2
timestamp 1666464484
transform -1 0 138880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__A3
timestamp 1666464484
transform 1 0 137312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__592__A1
timestamp 1666464484
transform 1 0 95760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__592__C
timestamp 1666464484
transform -1 0 100800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__593__A1
timestamp 1666464484
transform 1 0 95984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__A1
timestamp 1666464484
transform -1 0 130928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__A1
timestamp 1666464484
transform 1 0 100352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__A1
timestamp 1666464484
transform -1 0 100464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__A2
timestamp 1666464484
transform -1 0 95088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__B1
timestamp 1666464484
transform 1 0 93072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__C1
timestamp 1666464484
transform 1 0 101024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__C2
timestamp 1666464484
transform 1 0 98896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__597__A1
timestamp 1666464484
transform 1 0 92400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__597__A2
timestamp 1666464484
transform 1 0 93072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__A1
timestamp 1666464484
transform 1 0 100912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__A2
timestamp 1666464484
transform -1 0 99792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__A3
timestamp 1666464484
transform 1 0 99120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__598__A4
timestamp 1666464484
transform 1 0 100464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__A1
timestamp 1666464484
transform 1 0 100912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A1
timestamp 1666464484
transform -1 0 101248 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A2
timestamp 1666464484
transform -1 0 101696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__B1
timestamp 1666464484
transform -1 0 94304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__C1
timestamp 1666464484
transform -1 0 92848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__C2
timestamp 1666464484
transform -1 0 98336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__601__A1
timestamp 1666464484
transform -1 0 100016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A1
timestamp 1666464484
transform 1 0 101024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A2
timestamp 1666464484
transform 1 0 100464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__603__I
timestamp 1666464484
transform 1 0 100016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__A1
timestamp 1666464484
transform 1 0 95088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__A2
timestamp 1666464484
transform 1 0 93968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__A3
timestamp 1666464484
transform 1 0 94416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__I
timestamp 1666464484
transform -1 0 98448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__A1
timestamp 1666464484
transform 1 0 98672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__B
timestamp 1666464484
transform 1 0 100128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__607__A1
timestamp 1666464484
transform 1 0 102368 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__A1
timestamp 1666464484
transform -1 0 109648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__A2
timestamp 1666464484
transform -1 0 110880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__B2
timestamp 1666464484
transform 1 0 101920 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__609__B
timestamp 1666464484
transform 1 0 104384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__610__A1
timestamp 1666464484
transform 1 0 99792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__610__A2
timestamp 1666464484
transform 1 0 100240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__610__A3
timestamp 1666464484
transform 1 0 97664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__611__I
timestamp 1666464484
transform -1 0 94752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__A1
timestamp 1666464484
transform 1 0 96096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__A2
timestamp 1666464484
transform 1 0 94192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__B
timestamp 1666464484
transform 1 0 97776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__613__A1
timestamp 1666464484
transform 1 0 96656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__A1
timestamp 1666464484
transform -1 0 132384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__615__A1
timestamp 1666464484
transform -1 0 109984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__615__A2
timestamp 1666464484
transform -1 0 103040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__615__B2
timestamp 1666464484
transform 1 0 101472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__616__B
timestamp 1666464484
transform 1 0 100576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__I
timestamp 1666464484
transform 1 0 41888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__A1
timestamp 1666464484
transform 1 0 33488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__A2
timestamp 1666464484
transform 1 0 36288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__619__A1
timestamp 1666464484
transform -1 0 37072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__620__I
timestamp 1666464484
transform -1 0 63280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__621__I0
timestamp 1666464484
transform -1 0 61936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__I
timestamp 1666464484
transform -1 0 46144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__624__I
timestamp 1666464484
transform -1 0 23632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__625__I1
timestamp 1666464484
transform 1 0 15792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__625__S
timestamp 1666464484
transform -1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__I1
timestamp 1666464484
transform 1 0 18144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__S
timestamp 1666464484
transform 1 0 17696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__I1
timestamp 1666464484
transform 1 0 21952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__S
timestamp 1666464484
transform 1 0 21504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__I1
timestamp 1666464484
transform 1 0 24192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__S
timestamp 1666464484
transform 1 0 22848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__633__I
timestamp 1666464484
transform 1 0 30912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__I1
timestamp 1666464484
transform -1 0 26992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__636__A1
timestamp 1666464484
transform -1 0 37520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__636__A2
timestamp 1666464484
transform -1 0 39984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__637__A1
timestamp 1666464484
transform -1 0 36960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__I1
timestamp 1666464484
transform 1 0 27776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__640__I1
timestamp 1666464484
transform -1 0 29232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__642__A2
timestamp 1666464484
transform -1 0 31696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__643__A1
timestamp 1666464484
transform 1 0 36512 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__644__I1
timestamp 1666464484
transform -1 0 30688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__I
timestamp 1666464484
transform 1 0 32816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__I1
timestamp 1666464484
transform 1 0 35392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__649__I1
timestamp 1666464484
transform 1 0 35840 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__I
timestamp 1666464484
transform -1 0 44912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__A1
timestamp 1666464484
transform 1 0 42560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__A2
timestamp 1666464484
transform 1 0 43456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__653__A1
timestamp 1666464484
transform -1 0 42336 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__653__A2
timestamp 1666464484
transform -1 0 41664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__654__I
timestamp 1666464484
transform 1 0 43792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__A1
timestamp 1666464484
transform -1 0 51296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__A2
timestamp 1666464484
transform 1 0 50848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__A1
timestamp 1666464484
transform 1 0 54432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__A2
timestamp 1666464484
transform -1 0 52864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__I1
timestamp 1666464484
transform 1 0 39312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__I1
timestamp 1666464484
transform 1 0 41888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__661__I
timestamp 1666464484
transform -1 0 48832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__662__I1
timestamp 1666464484
transform -1 0 47264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__664__I1
timestamp 1666464484
transform 1 0 46368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__666__I1
timestamp 1666464484
transform 1 0 51072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__668__I1
timestamp 1666464484
transform 1 0 48720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__670__A2
timestamp 1666464484
transform -1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__671__A1
timestamp 1666464484
transform -1 0 44240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__671__A2
timestamp 1666464484
transform -1 0 42000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__A2
timestamp 1666464484
transform 1 0 50624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__A1
timestamp 1666464484
transform -1 0 52864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__A2
timestamp 1666464484
transform -1 0 51744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__I
timestamp 1666464484
transform 1 0 56336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__I1
timestamp 1666464484
transform 1 0 56000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__S
timestamp 1666464484
transform 1 0 56112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__I
timestamp 1666464484
transform 1 0 43008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__A2
timestamp 1666464484
transform 1 0 56784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__A1
timestamp 1666464484
transform -1 0 58464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__A2
timestamp 1666464484
transform -1 0 58016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__I1
timestamp 1666464484
transform -1 0 58016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__S
timestamp 1666464484
transform 1 0 57344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__I1
timestamp 1666464484
transform 1 0 59584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__S
timestamp 1666464484
transform 1 0 56672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__I0
timestamp 1666464484
transform 1 0 59136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__I1
timestamp 1666464484
transform 1 0 61936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__S
timestamp 1666464484
transform 1 0 59584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__A1
timestamp 1666464484
transform -1 0 59024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__A2
timestamp 1666464484
transform 1 0 59584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__A1
timestamp 1666464484
transform -1 0 62272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__A2
timestamp 1666464484
transform 1 0 59696 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__691__A1
timestamp 1666464484
transform -1 0 63504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__691__A2
timestamp 1666464484
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__692__CLK
timestamp 1666464484
transform -1 0 39200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__693__CLK
timestamp 1666464484
transform 1 0 58688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__694__CLK
timestamp 1666464484
transform 1 0 67088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__CLK
timestamp 1666464484
transform 1 0 68096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__696__CLK
timestamp 1666464484
transform 1 0 69216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__697__CLK
timestamp 1666464484
transform 1 0 65744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__CLK
timestamp 1666464484
transform 1 0 68544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__699__CLK
timestamp 1666464484
transform -1 0 72464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__700__CLK
timestamp 1666464484
transform -1 0 75600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__CLK
timestamp 1666464484
transform 1 0 76160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__702__CLK
timestamp 1666464484
transform 1 0 82992 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__703__CLK
timestamp 1666464484
transform 1 0 78848 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__704__CLK
timestamp 1666464484
transform 1 0 84448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__CLK
timestamp 1666464484
transform -1 0 88144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__706__CLK
timestamp 1666464484
transform 1 0 87584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__CLK
timestamp 1666464484
transform 1 0 81200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__CLK
timestamp 1666464484
transform 1 0 88928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__CLK
timestamp 1666464484
transform 1 0 102816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__CLK
timestamp 1666464484
transform -1 0 104608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__CLK
timestamp 1666464484
transform 1 0 107856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__D
timestamp 1666464484
transform 1 0 112672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__CLK
timestamp 1666464484
transform 1 0 108304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__D
timestamp 1666464484
transform 1 0 112784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__CLK
timestamp 1666464484
transform 1 0 108528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__D
timestamp 1666464484
transform -1 0 113232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__714__CLK
timestamp 1666464484
transform 1 0 107856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__CLK
timestamp 1666464484
transform 1 0 108304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__D
timestamp 1666464484
transform -1 0 112224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__CLK
timestamp 1666464484
transform 1 0 116032 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__717__CLK
timestamp 1666464484
transform 1 0 112784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__718__CLK
timestamp 1666464484
transform 1 0 101472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__CLK
timestamp 1666464484
transform 1 0 105504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__CLK
timestamp 1666464484
transform 1 0 93744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__721__CLK
timestamp 1666464484
transform 1 0 88480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__CLK
timestamp 1666464484
transform 1 0 98112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__CLK
timestamp 1666464484
transform 1 0 100352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__CLK
timestamp 1666464484
transform 1 0 96432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__725__CLK
timestamp 1666464484
transform 1 0 30688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__726__CLK
timestamp 1666464484
transform 1 0 62160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__727__CLK
timestamp 1666464484
transform -1 0 13888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__728__CLK
timestamp 1666464484
transform 1 0 17808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__CLK
timestamp 1666464484
transform 1 0 21504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__730__CLK
timestamp 1666464484
transform 1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__CLK
timestamp 1666464484
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__CLK
timestamp 1666464484
transform 1 0 38752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__733__CLK
timestamp 1666464484
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__CLK
timestamp 1666464484
transform 1 0 29008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__735__CLK
timestamp 1666464484
transform 1 0 35168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__736__CLK
timestamp 1666464484
transform 1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__CLK
timestamp 1666464484
transform 1 0 33936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__CLK
timestamp 1666464484
transform 1 0 32816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__739__CLK
timestamp 1666464484
transform 1 0 43120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__CLK
timestamp 1666464484
transform 1 0 45360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__741__CLK
timestamp 1666464484
transform 1 0 40880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__742__CLK
timestamp 1666464484
transform 1 0 41440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__743__CLK
timestamp 1666464484
transform -1 0 46704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__744__CLK
timestamp 1666464484
transform -1 0 46144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__746__CLK
timestamp 1666464484
transform -1 0 49952 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__747__CLK
timestamp 1666464484
transform 1 0 41664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__752__CLK
timestamp 1666464484
transform 1 0 56448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__753__CLK
timestamp 1666464484
transform 1 0 62832 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__754__CLK
timestamp 1666464484
transform 1 0 58240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__755__CLK
timestamp 1666464484
transform 1 0 63392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__756__CLK
timestamp 1666464484
transform 1 0 63728 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__799__I
timestamp 1666464484
transform 1 0 5152 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__800__I
timestamp 1666464484
transform 1 0 7952 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__801__I
timestamp 1666464484
transform 1 0 11088 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__802__I
timestamp 1666464484
transform 1 0 16016 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__803__I
timestamp 1666464484
transform 1 0 20832 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__804__I
timestamp 1666464484
transform 1 0 25536 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__805__I
timestamp 1666464484
transform 1 0 30240 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__806__I
timestamp 1666464484
transform 1 0 34608 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__807__I
timestamp 1666464484
transform 1 0 39648 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__808__I
timestamp 1666464484
transform 1 0 44352 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__809__I
timestamp 1666464484
transform 1 0 48720 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__810__I
timestamp 1666464484
transform 1 0 53760 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__811__I
timestamp 1666464484
transform 1 0 58128 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__812__I
timestamp 1666464484
transform 1 0 63168 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__813__I
timestamp 1666464484
transform 1 0 67872 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__814__I
timestamp 1666464484
transform 1 0 72576 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__815__I
timestamp 1666464484
transform 1 0 77280 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__816__I
timestamp 1666464484
transform 1 0 81648 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__817__I
timestamp 1666464484
transform 1 0 86688 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__818__I
timestamp 1666464484
transform 1 0 91392 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__819__I
timestamp 1666464484
transform 1 0 96432 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__820__I
timestamp 1666464484
transform 1 0 100800 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__821__I
timestamp 1666464484
transform 1 0 105392 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__822__I
timestamp 1666464484
transform 1 0 110432 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__823__I
timestamp 1666464484
transform 1 0 114912 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__824__I
timestamp 1666464484
transform 1 0 120288 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__825__I
timestamp 1666464484
transform 1 0 124208 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__826__I
timestamp 1666464484
transform 1 0 128912 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__827__I
timestamp 1666464484
transform 1 0 133728 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__828__I
timestamp 1666464484
transform 1 0 138432 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__829__I
timestamp 1666464484
transform 1 0 143136 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__830__I
timestamp 1666464484
transform 1 0 147840 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__831__I
timestamp 1666464484
transform 1 0 152096 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__832__I
timestamp 1666464484
transform 1 0 157248 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__833__I
timestamp 1666464484
transform 1 0 161952 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__834__I
timestamp 1666464484
transform 1 0 166656 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__835__I
timestamp 1666464484
transform 1 0 170016 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__836__I
timestamp 1666464484
transform 1 0 62608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__837__I
timestamp 1666464484
transform 1 0 64176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__838__I
timestamp 1666464484
transform 1 0 62496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__839__I
timestamp 1666464484
transform 1 0 64736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__840__I
timestamp 1666464484
transform 1 0 74144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__841__I
timestamp 1666464484
transform 1 0 74480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__842__I
timestamp 1666464484
transform 1 0 75824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__843__I
timestamp 1666464484
transform 1 0 75712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__844__I
timestamp 1666464484
transform 1 0 77392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__845__I
timestamp 1666464484
transform 1 0 80416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__846__I
timestamp 1666464484
transform 1 0 81424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__847__I
timestamp 1666464484
transform 1 0 82992 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__848__I
timestamp 1666464484
transform -1 0 81648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__849__I
timestamp 1666464484
transform 1 0 88480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__850__I
timestamp 1666464484
transform 1 0 90496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__851__I
timestamp 1666464484
transform -1 0 89264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__852__I
timestamp 1666464484
transform 1 0 93744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__853__I
timestamp 1666464484
transform 1 0 93520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__854__I
timestamp 1666464484
transform 1 0 100240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__855__I
timestamp 1666464484
transform 1 0 102816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__856__I
timestamp 1666464484
transform 1 0 101024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__857__I
timestamp 1666464484
transform 1 0 109872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__858__I
timestamp 1666464484
transform 1 0 114800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__859__I
timestamp 1666464484
transform 1 0 111216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__860__I
timestamp 1666464484
transform 1 0 106400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__861__I
timestamp 1666464484
transform 1 0 114352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__862__I
timestamp 1666464484
transform 1 0 114352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__863__I
timestamp 1666464484
transform 1 0 113232 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__864__I
timestamp 1666464484
transform 1 0 114128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__865__I
timestamp 1666464484
transform 1 0 114352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__866__I
timestamp 1666464484
transform 1 0 114800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__867__I
timestamp 1666464484
transform -1 0 117600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1666464484
transform 1 0 59248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1666464484
transform -1 0 55216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1666464484
transform 1 0 54992 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1666464484
transform 1 0 53648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1666464484
transform -1 0 48944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1666464484
transform -1 0 69664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1666464484
transform -1 0 68768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1666464484
transform 1 0 64176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1666464484
transform -1 0 69216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1666464484
transform 1 0 121520 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1666464484
transform -1 0 124432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1666464484
transform 1 0 125776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1666464484
transform -1 0 126224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1666464484
transform -1 0 128016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1666464484
transform 1 0 131376 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1666464484
transform -1 0 133056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1666464484
transform -1 0 133728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1666464484
transform 1 0 138880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1666464484
transform -1 0 137648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1666464484
transform 1 0 137648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1666464484
transform -1 0 141008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1666464484
transform 1 0 141904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1666464484
transform -1 0 141680 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1666464484
transform 1 0 144816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1666464484
transform -1 0 146384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1666464484
transform -1 0 147728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1666464484
transform -1 0 148848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1666464484
transform 1 0 151984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1666464484
transform -1 0 151312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1666464484
transform 1 0 154000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1666464484
transform -1 0 155456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1666464484
transform -1 0 155904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1666464484
transform -1 0 158480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1666464484
transform 1 0 160720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1666464484
transform -1 0 161168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1666464484
transform 1 0 164080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1666464484
transform 1 0 165760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1666464484
transform -1 0 167216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1666464484
transform -1 0 169456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1666464484
transform 1 0 170800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1666464484
transform 1 0 172480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1666464484
transform 1 0 123760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1666464484
transform 1 0 125440 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1666464484
transform 1 0 126448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1666464484
transform 1 0 127344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1666464484
transform -1 0 128912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1666464484
transform -1 0 132048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1666464484
transform 1 0 133168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1666464484
transform 1 0 135408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1666464484
transform -1 0 136752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1666464484
transform -1 0 138880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1666464484
transform -1 0 139776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1666464484
transform -1 0 140224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1666464484
transform 1 0 143024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1666464484
transform -1 0 143696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1666464484
transform -1 0 145488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1666464484
transform 1 0 147056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1666464484
transform 1 0 149968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1666464484
transform 1 0 150640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1666464484
transform 1 0 152768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1666464484
transform -1 0 152544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1666464484
transform -1 0 154672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1666464484
transform 1 0 156688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1666464484
transform 1 0 157696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1666464484
transform -1 0 159376 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1666464484
transform -1 0 161616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1666464484
transform 1 0 162736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1666464484
transform 1 0 164528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1666464484
transform -1 0 166432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1666464484
transform -1 0 168112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1666464484
transform -1 0 169008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1666464484
transform -1 0 171472 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1666464484
transform 1 0 173600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1666464484
transform -1 0 5936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1666464484
transform -1 0 7168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1666464484
transform -1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1666464484
transform -1 0 29680 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1666464484
transform -1 0 29680 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1666464484
transform -1 0 30128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1666464484
transform -1 0 31584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1666464484
transform -1 0 31696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1666464484
transform -1 0 36512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1666464484
transform -1 0 36736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1666464484
transform -1 0 36960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1666464484
transform -1 0 38864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1666464484
transform -1 0 44912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1666464484
transform -1 0 11872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1666464484
transform -1 0 44128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1666464484
transform -1 0 47264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1666464484
transform -1 0 47712 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1666464484
transform -1 0 41888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1666464484
transform -1 0 48160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1666464484
transform -1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1666464484
transform -1 0 55664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1666464484
transform -1 0 57568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1666464484
transform -1 0 57120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1666464484
transform 1 0 61264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1666464484
transform -1 0 14224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1666464484
transform -1 0 58464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1666464484
transform -1 0 64848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1666464484
transform -1 0 15008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1666464484
transform -1 0 17024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1666464484
transform -1 0 19936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1666464484
transform -1 0 22288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1666464484
transform -1 0 23968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1666464484
transform -1 0 23520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1666464484
transform -1 0 25424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1666464484
transform -1 0 10864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input100_I
timestamp 1666464484
transform -1 0 12768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input101_I
timestamp 1666464484
transform -1 0 15568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input102_I
timestamp 1666464484
transform -1 0 16464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input103_I
timestamp 1666464484
transform -1 0 8064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input104_I
timestamp 1666464484
transform 1 0 9632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output142_I
timestamp 1666464484
transform 1 0 6608 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output143_I
timestamp 1666464484
transform 1 0 55104 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output144_I
timestamp 1666464484
transform 1 0 58352 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output145_I
timestamp 1666464484
transform 1 0 62832 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output146_I
timestamp 1666464484
transform 1 0 67536 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output147_I
timestamp 1666464484
transform 1 0 72240 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output148_I
timestamp 1666464484
transform 1 0 78624 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output149_I
timestamp 1666464484
transform 1 0 81872 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output150_I
timestamp 1666464484
transform 1 0 86352 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output151_I
timestamp 1666464484
transform 1 0 91056 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output152_I
timestamp 1666464484
transform -1 0 95984 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output153_I
timestamp 1666464484
transform 1 0 11312 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output154_I
timestamp 1666464484
transform 1 0 102144 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output155_I
timestamp 1666464484
transform 1 0 105392 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output156_I
timestamp 1666464484
transform -1 0 110096 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output157_I
timestamp 1666464484
transform 1 0 113008 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output158_I
timestamp 1666464484
transform -1 0 117264 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output159_I
timestamp 1666464484
transform 1 0 122528 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output160_I
timestamp 1666464484
transform 1 0 126896 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output161_I
timestamp 1666464484
transform -1 0 131376 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output162_I
timestamp 1666464484
transform 1 0 136864 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output163_I
timestamp 1666464484
transform -1 0 140784 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output164_I
timestamp 1666464484
transform 1 0 15792 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output165_I
timestamp 1666464484
transform 1 0 146048 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output166_I
timestamp 1666464484
transform 1 0 150416 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output167_I
timestamp 1666464484
transform 1 0 20496 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output168_I
timestamp 1666464484
transform 1 0 25200 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output169_I
timestamp 1666464484
transform 1 0 31584 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output170_I
timestamp 1666464484
transform 1 0 34832 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output171_I
timestamp 1666464484
transform 1 0 39312 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output172_I
timestamp 1666464484
transform 1 0 44016 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output173_I
timestamp 1666464484
transform 1 0 48720 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output206_I
timestamp 1666464484
transform -1 0 6944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output207_I
timestamp 1666464484
transform 1 0 11200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output212_I
timestamp 1666464484
transform -1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output213_I
timestamp 1666464484
transform -1 0 32144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output218_I
timestamp 1666464484
transform 1 0 11984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output227_I
timestamp 1666464484
transform 1 0 60256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output236_I
timestamp 1666464484
transform -1 0 21952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41
timestamp 1666464484
transform 1 0 5936 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1666464484
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72
timestamp 1666464484
transform 1 0 9408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88
timestamp 1666464484
transform 1 0 11200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1666464484
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107
timestamp 1666464484
transform 1 0 13328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109
timestamp 1666464484
transform 1 0 13552 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112
timestamp 1666464484
transform 1 0 13888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120
timestamp 1666464484
transform 1 0 14784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_136 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 16576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1666464484
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_157
timestamp 1666464484
transform 1 0 18928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_159
timestamp 1666464484
transform 1 0 19152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1666464484
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1666464484
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_193
timestamp 1666464484
transform 1 0 22960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1666464484
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1666464484
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_219
timestamp 1666464484
transform 1 0 25872 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_236
timestamp 1666464484
transform 1 0 27776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1666464484
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_247
timestamp 1666464484
transform 1 0 29008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_255
timestamp 1666464484
transform 1 0 29904 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_272
timestamp 1666464484
transform 1 0 31808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_276
timestamp 1666464484
transform 1 0 32256 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1666464484
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1666464484
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_297
timestamp 1666464484
transform 1 0 34608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_299
timestamp 1666464484
transform 1 0 34832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1666464484
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317
timestamp 1666464484
transform 1 0 36848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_333
timestamp 1666464484
transform 1 0 38640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_352
timestamp 1666464484
transform 1 0 40768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_368
timestamp 1666464484
transform 1 0 42560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1666464484
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_387
timestamp 1666464484
transform 1 0 44688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_403
timestamp 1666464484
transform 1 0 46480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_422
timestamp 1666464484
transform 1 0 48608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_424
timestamp 1666464484
transform 1 0 48832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1666464484
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_457
timestamp 1666464484
transform 1 0 52528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_473
timestamp 1666464484
transform 1 0 54320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1666464484
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_492
timestamp 1666464484
transform 1 0 56448 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_508
timestamp 1666464484
transform 1 0 58240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_524
timestamp 1666464484
transform 1 0 60032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_527
timestamp 1666464484
transform 1 0 60368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_543
timestamp 1666464484
transform 1 0 62160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1666464484
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_562
timestamp 1666464484
transform 1 0 64288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_564
timestamp 1666464484
transform 1 0 64512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_567
timestamp 1666464484
transform 1 0 64848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_575
timestamp 1666464484
transform 1 0 65744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_591
timestamp 1666464484
transform 1 0 67536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1666464484
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_612
timestamp 1666464484
transform 1 0 69888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_614
timestamp 1666464484
transform 1 0 70112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1666464484
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_632
timestamp 1666464484
transform 1 0 72128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_648
timestamp 1666464484
transform 1 0 73920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1666464484
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_667
timestamp 1666464484
transform 1 0 76048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_669
timestamp 1666464484
transform 1 0 76272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_672
timestamp 1666464484
transform 1 0 76608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_680
timestamp 1666464484
transform 1 0 77504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_696
timestamp 1666464484
transform 1 0 79296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_702
timestamp 1666464484
transform 1 0 79968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_718
timestamp 1666464484
transform 1 0 81760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_734
timestamp 1666464484
transform 1 0 83552 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_737
timestamp 1666464484
transform 1 0 83888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_753
timestamp 1666464484
transform 1 0 85680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_769
timestamp 1666464484
transform 1 0 87472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_772
timestamp 1666464484
transform 1 0 87808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_774
timestamp 1666464484
transform 1 0 88032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_777
timestamp 1666464484
transform 1 0 88368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_781
timestamp 1666464484
transform 1 0 88816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_785
timestamp 1666464484
transform 1 0 89264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_801
timestamp 1666464484
transform 1 0 91056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_807
timestamp 1666464484
transform 1 0 91728 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_822
timestamp 1666464484
transform 1 0 93408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_838
timestamp 1666464484
transform 1 0 95200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_842
timestamp 1666464484
transform 1 0 95648 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_845
timestamp 1666464484
transform 1 0 95984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_861
timestamp 1666464484
transform 1 0 97776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_869
timestamp 1666464484
transform 1 0 98672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_873
timestamp 1666464484
transform 1 0 99120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_877
timestamp 1666464484
transform 1 0 99568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_892
timestamp 1666464484
transform 1 0 101248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_908
timestamp 1666464484
transform 1 0 103040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_912
timestamp 1666464484
transform 1 0 103488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_927
timestamp 1666464484
transform 1 0 105168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_943
timestamp 1666464484
transform 1 0 106960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_947
timestamp 1666464484
transform 1 0 107408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_950
timestamp 1666464484
transform 1 0 107744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_966
timestamp 1666464484
transform 1 0 109536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_970
timestamp 1666464484
transform 1 0 109984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_974
timestamp 1666464484
transform 1 0 110432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_978
timestamp 1666464484
transform 1 0 110880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1666464484
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_997
timestamp 1666464484
transform 1 0 113008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1013
timestamp 1666464484
transform 1 0 114800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1017
timestamp 1666464484
transform 1 0 115248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1032
timestamp 1666464484
transform 1 0 116928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1048
timestamp 1666464484
transform 1 0 118720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1052
timestamp 1666464484
transform 1 0 119168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1067
timestamp 1666464484
transform 1 0 120848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1078
timestamp 1666464484
transform 1 0 122080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1084
timestamp 1666464484
transform 1 0 122752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1087
timestamp 1666464484
transform 1 0 123088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1094
timestamp 1666464484
transform 1 0 123872 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1102
timestamp 1666464484
transform 1 0 124768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1110
timestamp 1666464484
transform 1 0 125664 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1118
timestamp 1666464484
transform 1 0 126560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1122
timestamp 1666464484
transform 1 0 127008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1129
timestamp 1666464484
transform 1 0 127792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1137
timestamp 1666464484
transform 1 0 128688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1145
timestamp 1666464484
transform 1 0 129584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1153
timestamp 1666464484
transform 1 0 130480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1157
timestamp 1666464484
transform 1 0 130928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1164
timestamp 1666464484
transform 1 0 131712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1172
timestamp 1666464484
transform 1 0 132608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1180
timestamp 1666464484
transform 1 0 133504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1188
timestamp 1666464484
transform 1 0 134400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1192
timestamp 1666464484
transform 1 0 134848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1199
timestamp 1666464484
transform 1 0 135632 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1207
timestamp 1666464484
transform 1 0 136528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1215
timestamp 1666464484
transform 1 0 137424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1223
timestamp 1666464484
transform 1 0 138320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1227
timestamp 1666464484
transform 1 0 138768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1234
timestamp 1666464484
transform 1 0 139552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1242
timestamp 1666464484
transform 1 0 140448 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1250
timestamp 1666464484
transform 1 0 141344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1258
timestamp 1666464484
transform 1 0 142240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1262
timestamp 1666464484
transform 1 0 142688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1269
timestamp 1666464484
transform 1 0 143472 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1277
timestamp 1666464484
transform 1 0 144368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1285
timestamp 1666464484
transform 1 0 145264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1293
timestamp 1666464484
transform 1 0 146160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1297
timestamp 1666464484
transform 1 0 146608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1304
timestamp 1666464484
transform 1 0 147392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1312
timestamp 1666464484
transform 1 0 148288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1320
timestamp 1666464484
transform 1 0 149184 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1328
timestamp 1666464484
transform 1 0 150080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1332
timestamp 1666464484
transform 1 0 150528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1339
timestamp 1666464484
transform 1 0 151312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1347
timestamp 1666464484
transform 1 0 152208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1355
timestamp 1666464484
transform 1 0 153104 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1363
timestamp 1666464484
transform 1 0 154000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1367
timestamp 1666464484
transform 1 0 154448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1374
timestamp 1666464484
transform 1 0 155232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1382
timestamp 1666464484
transform 1 0 156128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1390
timestamp 1666464484
transform 1 0 157024 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1398
timestamp 1666464484
transform 1 0 157920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1402
timestamp 1666464484
transform 1 0 158368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1409
timestamp 1666464484
transform 1 0 159152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1417
timestamp 1666464484
transform 1 0 160048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1425
timestamp 1666464484
transform 1 0 160944 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1433
timestamp 1666464484
transform 1 0 161840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1437
timestamp 1666464484
transform 1 0 162288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1444
timestamp 1666464484
transform 1 0 163072 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1452
timestamp 1666464484
transform 1 0 163968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1460
timestamp 1666464484
transform 1 0 164864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1468
timestamp 1666464484
transform 1 0 165760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1472
timestamp 1666464484
transform 1 0 166208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1479
timestamp 1666464484
transform 1 0 166992 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1487
timestamp 1666464484
transform 1 0 167888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1495
timestamp 1666464484
transform 1 0 168784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1503
timestamp 1666464484
transform 1 0 169680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1507
timestamp 1666464484
transform 1 0 170128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1514
timestamp 1666464484
transform 1 0 170912 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1522
timestamp 1666464484
transform 1 0 171808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1530
timestamp 1666464484
transform 1 0 172704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1538
timestamp 1666464484
transform 1 0 173600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1542
timestamp 1666464484
transform 1 0 174048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1547
timestamp 1666464484
transform 1 0 174608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1553 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 175280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1569
timestamp 1666464484
transform 1 0 177072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1573
timestamp 1666464484
transform 1 0 177520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1577
timestamp 1666464484
transform 1 0 177968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_2
timestamp 1666464484
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_34 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5152 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_42
timestamp 1666464484
transform 1 0 6048 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_46
timestamp 1666464484
transform 1 0 6496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_50
timestamp 1666464484
transform 1 0 6944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_66
timestamp 1666464484
transform 1 0 8736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1666464484
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_73
timestamp 1666464484
transform 1 0 9520 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_83
timestamp 1666464484
transform 1 0 10640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_85
timestamp 1666464484
transform 1 0 10864 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_92
timestamp 1666464484
transform 1 0 11648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_123
timestamp 1666464484
transform 1 0 15120 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_133
timestamp 1666464484
transform 1 0 16240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1666464484
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_144
timestamp 1666464484
transform 1 0 17472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_146
timestamp 1666464484
transform 1 0 17696 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_149
timestamp 1666464484
transform 1 0 18032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_157
timestamp 1666464484
transform 1 0 18928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_188
timestamp 1666464484
transform 1 0 22400 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_196
timestamp 1666464484
transform 1 0 23296 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1666464484
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1666464484
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_222
timestamp 1666464484
transform 1 0 26208 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_239
timestamp 1666464484
transform 1 0 28112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_245
timestamp 1666464484
transform 1 0 28784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_276
timestamp 1666464484
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_280
timestamp 1666464484
transform 1 0 32704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1666464484
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1666464484
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_289
timestamp 1666464484
transform 1 0 33712 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_305
timestamp 1666464484
transform 1 0 35504 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_336
timestamp 1666464484
transform 1 0 38976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_343
timestamp 1666464484
transform 1 0 39760 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1666464484
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_357
timestamp 1666464484
transform 1 0 41328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_359
timestamp 1666464484
transform 1 0 41552 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_362
timestamp 1666464484
transform 1 0 41888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_375
timestamp 1666464484
transform 1 0 43344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_391
timestamp 1666464484
transform 1 0 45136 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_422
timestamp 1666464484
transform 1 0 48608 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1666464484
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_479
timestamp 1666464484
transform 1 0 54992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_495
timestamp 1666464484
transform 1 0 56784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1666464484
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_506
timestamp 1666464484
transform 1 0 58016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_537
timestamp 1666464484
transform 1 0 61488 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_541
timestamp 1666464484
transform 1 0 61936 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_549
timestamp 1666464484
transform 1 0 62832 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_557
timestamp 1666464484
transform 1 0 63728 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_565
timestamp 1666464484
transform 1 0 64624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1666464484
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1666464484
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_585
timestamp 1666464484
transform 1 0 66864 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_600
timestamp 1666464484
transform 1 0 68544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_604
timestamp 1666464484
transform 1 0 68992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_620
timestamp 1666464484
transform 1 0 70784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_636
timestamp 1666464484
transform 1 0 72576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1666464484
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1666464484
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_656
timestamp 1666464484
transform 1 0 74816 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_658
timestamp 1666464484
transform 1 0 75040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_665
timestamp 1666464484
transform 1 0 75824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_681
timestamp 1666464484
transform 1 0 77616 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_685
timestamp 1666464484
transform 1 0 78064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_693
timestamp 1666464484
transform 1 0 78960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_709
timestamp 1666464484
transform 1 0 80752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_712
timestamp 1666464484
transform 1 0 81088 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_714
timestamp 1666464484
transform 1 0 81312 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_717
timestamp 1666464484
transform 1 0 81648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_725
timestamp 1666464484
transform 1 0 82544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_738
timestamp 1666464484
transform 1 0 84000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_754
timestamp 1666464484
transform 1 0 85792 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_764
timestamp 1666464484
transform 1 0 86912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_780
timestamp 1666464484
transform 1 0 88704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_783
timestamp 1666464484
transform 1 0 89040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_788
timestamp 1666464484
transform 1 0 89600 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_804
timestamp 1666464484
transform 1 0 91392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_812
timestamp 1666464484
transform 1 0 92288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_814
timestamp 1666464484
transform 1 0 92512 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_823
timestamp 1666464484
transform 1 0 93520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_827
timestamp 1666464484
transform 1 0 93968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_831
timestamp 1666464484
transform 1 0 94416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_846
timestamp 1666464484
transform 1 0 96096 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_850
timestamp 1666464484
transform 1 0 96544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_854
timestamp 1666464484
transform 1 0 96992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_860
timestamp 1666464484
transform 1 0 97664 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_876
timestamp 1666464484
transform 1 0 99456 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_887
timestamp 1666464484
transform 1 0 100688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_893
timestamp 1666464484
transform 1 0 101360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_904
timestamp 1666464484
transform 1 0 102592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_912
timestamp 1666464484
transform 1 0 103488 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_922
timestamp 1666464484
transform 1 0 104608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_925
timestamp 1666464484
transform 1 0 104944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_927
timestamp 1666464484
transform 1 0 105168 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_935
timestamp 1666464484
transform 1 0 106064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_951
timestamp 1666464484
transform 1 0 107856 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_967
timestamp 1666464484
transform 1 0 109648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_983
timestamp 1666464484
transform 1 0 111440 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_993
timestamp 1666464484
transform 1 0 112560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_996
timestamp 1666464484
transform 1 0 112896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1011
timestamp 1666464484
transform 1 0 114576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1015
timestamp 1666464484
transform 1 0 115024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1017
timestamp 1666464484
transform 1 0 115248 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1032
timestamp 1666464484
transform 1 0 116928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1048
timestamp 1666464484
transform 1 0 118720 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1052
timestamp 1666464484
transform 1 0 119168 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1064
timestamp 1666464484
transform 1 0 120512 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1067
timestamp 1666464484
transform 1 0 120848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1082
timestamp 1666464484
transform 1 0 122528 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1086
timestamp 1666464484
transform 1 0 122976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1088
timestamp 1666464484
transform 1 0 123200 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1097
timestamp 1666464484
transform 1 0 124208 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1105
timestamp 1666464484
transform 1 0 125104 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1113
timestamp 1666464484
transform 1 0 126000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1121
timestamp 1666464484
transform 1 0 126896 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1125
timestamp 1666464484
transform 1 0 127344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1133
timestamp 1666464484
transform 1 0 128240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1135
timestamp 1666464484
transform 1 0 128464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1138
timestamp 1666464484
transform 1 0 128800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1145
timestamp 1666464484
transform 1 0 129584 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1153
timestamp 1666464484
transform 1 0 130480 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1161
timestamp 1666464484
transform 1 0 131376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1169
timestamp 1666464484
transform 1 0 132272 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1177
timestamp 1666464484
transform 1 0 133168 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1185
timestamp 1666464484
transform 1 0 134064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1193
timestamp 1666464484
transform 1 0 134960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1201
timestamp 1666464484
transform 1 0 135856 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1205
timestamp 1666464484
transform 1 0 136304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1209
timestamp 1666464484
transform 1 0 136752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1218
timestamp 1666464484
transform 1 0 137760 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1230
timestamp 1666464484
transform 1 0 139104 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1238
timestamp 1666464484
transform 1 0 140000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1246
timestamp 1666464484
transform 1 0 140896 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1250
timestamp 1666464484
transform 1 0 141344 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1261
timestamp 1666464484
transform 1 0 142576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1271
timestamp 1666464484
transform 1 0 143696 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1277
timestamp 1666464484
transform 1 0 144368 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1280
timestamp 1666464484
transform 1 0 144704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1289
timestamp 1666464484
transform 1 0 145712 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1297
timestamp 1666464484
transform 1 0 146608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1305
timestamp 1666464484
transform 1 0 147504 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1313
timestamp 1666464484
transform 1 0 148400 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1321
timestamp 1666464484
transform 1 0 149296 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1329
timestamp 1666464484
transform 1 0 150192 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1335
timestamp 1666464484
transform 1 0 150864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1343
timestamp 1666464484
transform 1 0 151760 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1347
timestamp 1666464484
transform 1 0 152208 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1351
timestamp 1666464484
transform 1 0 152656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1354
timestamp 1666464484
transform 1 0 152992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1356
timestamp 1666464484
transform 1 0 153216 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1361
timestamp 1666464484
transform 1 0 153776 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1365
timestamp 1666464484
transform 1 0 154224 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1369
timestamp 1666464484
transform 1 0 154672 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1371
timestamp 1666464484
transform 1 0 154896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1376
timestamp 1666464484
transform 1 0 155456 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1380
timestamp 1666464484
transform 1 0 155904 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1388
timestamp 1666464484
transform 1 0 156800 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1394
timestamp 1666464484
transform 1 0 157472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1398
timestamp 1666464484
transform 1 0 157920 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1400
timestamp 1666464484
transform 1 0 158144 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1405
timestamp 1666464484
transform 1 0 158704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1411
timestamp 1666464484
transform 1 0 159376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1419
timestamp 1666464484
transform 1 0 160272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1422
timestamp 1666464484
transform 1 0 160608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1425
timestamp 1666464484
transform 1 0 160944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1433
timestamp 1666464484
transform 1 0 161840 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1439
timestamp 1666464484
transform 1 0 162512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1443
timestamp 1666464484
transform 1 0 162960 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1451
timestamp 1666464484
transform 1 0 163856 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1455
timestamp 1666464484
transform 1 0 164304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1459
timestamp 1666464484
transform 1 0 164752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1461
timestamp 1666464484
transform 1 0 164976 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1466
timestamp 1666464484
transform 1 0 165536 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1470
timestamp 1666464484
transform 1 0 165984 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1474
timestamp 1666464484
transform 1 0 166432 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1476
timestamp 1666464484
transform 1 0 166656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1481
timestamp 1666464484
transform 1 0 167216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1485
timestamp 1666464484
transform 1 0 167664 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1490
timestamp 1666464484
transform 1 0 168224 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1493
timestamp 1666464484
transform 1 0 168560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1503
timestamp 1666464484
transform 1 0 169680 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1511
timestamp 1666464484
transform 1 0 170576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1515
timestamp 1666464484
transform 1 0 171024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1519
timestamp 1666464484
transform 1 0 171472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1521
timestamp 1666464484
transform 1 0 171696 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1526
timestamp 1666464484
transform 1 0 172256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1530
timestamp 1666464484
transform 1 0 172704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1536
timestamp 1666464484
transform 1 0 173376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1540
timestamp 1666464484
transform 1 0 173824 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1556
timestamp 1666464484
transform 1 0 175616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1560
timestamp 1666464484
transform 1 0 176064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1564
timestamp 1666464484
transform 1 0 176512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1580
timestamp 1666464484
transform 1 0 178304 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1666464484
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1666464484
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_37
timestamp 1666464484
transform 1 0 5488 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_45
timestamp 1666464484
transform 1 0 6384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_49
timestamp 1666464484
transform 1 0 6832 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_52
timestamp 1666464484
transform 1 0 7168 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_60
timestamp 1666464484
transform 1 0 8064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_70
timestamp 1666464484
transform 1 0 9184 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_78
timestamp 1666464484
transform 1 0 10080 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_82
timestamp 1666464484
transform 1 0 10528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_85
timestamp 1666464484
transform 1 0 10864 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_93
timestamp 1666464484
transform 1 0 11760 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_97
timestamp 1666464484
transform 1 0 12208 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1666464484
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1666464484
transform 1 0 13440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_111
timestamp 1666464484
transform 1 0 13776 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_128
timestamp 1666464484
transform 1 0 15680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_159
timestamp 1666464484
transform 1 0 19152 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_161
timestamp 1666464484
transform 1 0 19376 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_179
timestamp 1666464484
transform 1 0 21392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_181
timestamp 1666464484
transform 1 0 21616 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_184
timestamp 1666464484
transform 1 0 21952 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_200
timestamp 1666464484
transform 1 0 23744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_231
timestamp 1666464484
transform 1 0 27216 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1666464484
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_250
timestamp 1666464484
transform 1 0 29344 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_260
timestamp 1666464484
transform 1 0 30464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_264
timestamp 1666464484
transform 1 0 30912 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_280
timestamp 1666464484
transform 1 0 32704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_311
timestamp 1666464484
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_315
timestamp 1666464484
transform 1 0 36624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1666464484
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1666464484
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_330
timestamp 1666464484
transform 1 0 38304 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_338
timestamp 1666464484
transform 1 0 39200 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_346
timestamp 1666464484
transform 1 0 40096 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_377
timestamp 1666464484
transform 1 0 43568 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_381
timestamp 1666464484
transform 1 0 44016 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1666464484
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1666464484
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_395
timestamp 1666464484
transform 1 0 45584 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_403
timestamp 1666464484
transform 1 0 46480 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_419
timestamp 1666464484
transform 1 0 48272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_429
timestamp 1666464484
transform 1 0 49392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1666464484
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_463
timestamp 1666464484
transform 1 0 53200 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_496
timestamp 1666464484
transform 1 0 56896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_500
timestamp 1666464484
transform 1 0 57344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1666464484
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_550
timestamp 1666464484
transform 1 0 62944 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_554
timestamp 1666464484
transform 1 0 63392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_557
timestamp 1666464484
transform 1 0 63728 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_565
timestamp 1666464484
transform 1 0 64624 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_573
timestamp 1666464484
transform 1 0 65520 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_587
timestamp 1666464484
transform 1 0 67088 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1666464484
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1666464484
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_617
timestamp 1666464484
transform 1 0 70448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_626
timestamp 1666464484
transform 1 0 71456 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_628
timestamp 1666464484
transform 1 0 71680 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_661
timestamp 1666464484
transform 1 0 75376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_665
timestamp 1666464484
transform 1 0 75824 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1666464484
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_676
timestamp 1666464484
transform 1 0 77056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_691
timestamp 1666464484
transform 1 0 78736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_699
timestamp 1666464484
transform 1 0 79632 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_707
timestamp 1666464484
transform 1 0 80528 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_715
timestamp 1666464484
transform 1 0 81424 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_723
timestamp 1666464484
transform 1 0 82320 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_725
timestamp 1666464484
transform 1 0 82544 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_728
timestamp 1666464484
transform 1 0 82880 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1666464484
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_747
timestamp 1666464484
transform 1 0 85008 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_749
timestamp 1666464484
transform 1 0 85232 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_756
timestamp 1666464484
transform 1 0 86016 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_772
timestamp 1666464484
transform 1 0 87808 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_774
timestamp 1666464484
transform 1 0 88032 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_777
timestamp 1666464484
transform 1 0 88368 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_791
timestamp 1666464484
transform 1 0 89936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_807
timestamp 1666464484
transform 1 0 91728 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1666464484
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_818
timestamp 1666464484
transform 1 0 92960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_825
timestamp 1666464484
transform 1 0 93744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_833
timestamp 1666464484
transform 1 0 94640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_841
timestamp 1666464484
transform 1 0 95536 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_849
timestamp 1666464484
transform 1 0 96432 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_865
timestamp 1666464484
transform 1 0 98224 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_881
timestamp 1666464484
transform 1 0 100016 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_885
timestamp 1666464484
transform 1 0 100464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_889
timestamp 1666464484
transform 1 0 100912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_892
timestamp 1666464484
transform 1 0 101248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_905
timestamp 1666464484
transform 1 0 102704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_925
timestamp 1666464484
transform 1 0 104944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_941
timestamp 1666464484
transform 1 0 106736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_943
timestamp 1666464484
transform 1 0 106960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_957
timestamp 1666464484
transform 1 0 108528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_960
timestamp 1666464484
transform 1 0 108864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_967
timestamp 1666464484
transform 1 0 109648 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_977
timestamp 1666464484
transform 1 0 110768 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_985
timestamp 1666464484
transform 1 0 111664 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_999
timestamp 1666464484
transform 1 0 113232 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1013
timestamp 1666464484
transform 1 0 114800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1021
timestamp 1666464484
transform 1 0 115696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1025
timestamp 1666464484
transform 1 0 116144 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1031
timestamp 1666464484
transform 1 0 116816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1038
timestamp 1666464484
transform 1 0 117600 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1042
timestamp 1666464484
transform 1 0 118048 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1049
timestamp 1666464484
transform 1 0 118832 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1062
timestamp 1666464484
transform 1 0 120288 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1078
timestamp 1666464484
transform 1 0 122080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1084
timestamp 1666464484
transform 1 0 122752 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1098
timestamp 1666464484
transform 1 0 124320 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1102
timestamp 1666464484
transform 1 0 124768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1115
timestamp 1666464484
transform 1 0 126224 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1121
timestamp 1666464484
transform 1 0 126896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1123
timestamp 1666464484
transform 1 0 127120 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1136
timestamp 1666464484
transform 1 0 128576 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1144
timestamp 1666464484
transform 1 0 129472 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1150
timestamp 1666464484
transform 1 0 130144 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1160
timestamp 1666464484
transform 1 0 131264 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1168
timestamp 1666464484
transform 1 0 132160 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1170
timestamp 1666464484
transform 1 0 132384 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1173
timestamp 1666464484
transform 1 0 132720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1184
timestamp 1666464484
transform 1 0 133952 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1192
timestamp 1666464484
transform 1 0 134848 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1204
timestamp 1666464484
transform 1 0 136192 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1216
timestamp 1666464484
transform 1 0 137536 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1227
timestamp 1666464484
transform 1 0 138768 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1235
timestamp 1666464484
transform 1 0 139664 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1241
timestamp 1666464484
transform 1 0 140336 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1244
timestamp 1666464484
transform 1 0 140672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1251
timestamp 1666464484
transform 1 0 141456 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1259
timestamp 1666464484
transform 1 0 142352 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1261
timestamp 1666464484
transform 1 0 142576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1270
timestamp 1666464484
transform 1 0 143584 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1278
timestamp 1666464484
transform 1 0 144480 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1280
timestamp 1666464484
transform 1 0 144704 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1287
timestamp 1666464484
transform 1 0 145488 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1295
timestamp 1666464484
transform 1 0 146384 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1303
timestamp 1666464484
transform 1 0 147280 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1311
timestamp 1666464484
transform 1 0 148176 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1315
timestamp 1666464484
transform 1 0 148624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1322
timestamp 1666464484
transform 1 0 149408 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1326
timestamp 1666464484
transform 1 0 149856 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1331
timestamp 1666464484
transform 1 0 150416 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1335
timestamp 1666464484
transform 1 0 150864 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1339
timestamp 1666464484
transform 1 0 151312 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1341
timestamp 1666464484
transform 1 0 151536 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1346
timestamp 1666464484
transform 1 0 152096 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1350
timestamp 1666464484
transform 1 0 152544 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1366
timestamp 1666464484
transform 1 0 154336 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1376
timestamp 1666464484
transform 1 0 155456 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1386
timestamp 1666464484
transform 1 0 156576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1389
timestamp 1666464484
transform 1 0 156912 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1397
timestamp 1666464484
transform 1 0 157808 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1403
timestamp 1666464484
transform 1 0 158480 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1407
timestamp 1666464484
transform 1 0 158928 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1411
timestamp 1666464484
transform 1 0 159376 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1419
timestamp 1666464484
transform 1 0 160272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1423
timestamp 1666464484
transform 1 0 160720 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1427
timestamp 1666464484
transform 1 0 161168 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1431
timestamp 1666464484
transform 1 0 161616 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1447
timestamp 1666464484
transform 1 0 163408 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1457
timestamp 1666464484
transform 1 0 164528 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1473
timestamp 1666464484
transform 1 0 166320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1477
timestamp 1666464484
transform 1 0 166768 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1481
timestamp 1666464484
transform 1 0 167216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1485
timestamp 1666464484
transform 1 0 167664 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1489
timestamp 1666464484
transform 1 0 168112 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1493
timestamp 1666464484
transform 1 0 168560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1497
timestamp 1666464484
transform 1 0 169008 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1501
timestamp 1666464484
transform 1 0 169456 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1517
timestamp 1666464484
transform 1 0 171248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1525
timestamp 1666464484
transform 1 0 172144 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_1528
timestamp 1666464484
transform 1 0 172480 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1560
timestamp 1666464484
transform 1 0 176064 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1576
timestamp 1666464484
transform 1 0 177856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1580
timestamp 1666464484
transform 1 0 178304 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_2
timestamp 1666464484
transform 1 0 1568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_34
timestamp 1666464484
transform 1 0 5152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_50
timestamp 1666464484
transform 1 0 6944 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_60
timestamp 1666464484
transform 1 0 8064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_68
timestamp 1666464484
transform 1 0 8960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1666464484
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1666464484
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_76
timestamp 1666464484
transform 1 0 9856 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_84
timestamp 1666464484
transform 1 0 10752 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_90
timestamp 1666464484
transform 1 0 11424 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_94
timestamp 1666464484
transform 1 0 11872 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_98
timestamp 1666464484
transform 1 0 12320 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_102
timestamp 1666464484
transform 1 0 12768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_110
timestamp 1666464484
transform 1 0 13664 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_118
timestamp 1666464484
transform 1 0 14560 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_125
timestamp 1666464484
transform 1 0 15344 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_133
timestamp 1666464484
transform 1 0 16240 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_140
timestamp 1666464484
transform 1 0 17024 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1666464484
transform 1 0 17472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_160
timestamp 1666464484
transform 1 0 19264 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_166
timestamp 1666464484
transform 1 0 19936 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_174
timestamp 1666464484
transform 1 0 20832 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_182
timestamp 1666464484
transform 1 0 21728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_186
timestamp 1666464484
transform 1 0 22176 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_193
timestamp 1666464484
transform 1 0 22960 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_199
timestamp 1666464484
transform 1 0 23632 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_201
timestamp 1666464484
transform 1 0 23856 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_208
timestamp 1666464484
transform 1 0 24640 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1666464484
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1666464484
transform 1 0 25424 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_245
timestamp 1666464484
transform 1 0 28784 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_249
timestamp 1666464484
transform 1 0 29232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_251
timestamp 1666464484
transform 1 0 29456 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_266
timestamp 1666464484
transform 1 0 31136 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_268
timestamp 1666464484
transform 1 0 31360 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_271
timestamp 1666464484
transform 1 0 31696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_275
timestamp 1666464484
transform 1 0 32144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1666464484
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_286
timestamp 1666464484
transform 1 0 33376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_288
timestamp 1666464484
transform 1 0 33600 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_295
timestamp 1666464484
transform 1 0 34384 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_303
timestamp 1666464484
transform 1 0 35280 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_334
timestamp 1666464484
transform 1 0 38752 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_342
timestamp 1666464484
transform 1 0 39648 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_346
timestamp 1666464484
transform 1 0 40096 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1666464484
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_357
timestamp 1666464484
transform 1 0 41328 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_363
timestamp 1666464484
transform 1 0 42000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_376
timestamp 1666464484
transform 1 0 43456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_380
timestamp 1666464484
transform 1 0 43904 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_383
timestamp 1666464484
transform 1 0 44240 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_393
timestamp 1666464484
transform 1 0 45360 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_397
timestamp 1666464484
transform 1 0 45808 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_400
timestamp 1666464484
transform 1 0 46144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_408
timestamp 1666464484
transform 1 0 47040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_418
timestamp 1666464484
transform 1 0 48160 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_422
timestamp 1666464484
transform 1 0 48608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1666464484
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1666464484
transform 1 0 49280 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_479
timestamp 1666464484
transform 1 0 54992 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1666464484
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1666464484
transform 1 0 57232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_508
timestamp 1666464484
transform 1 0 58240 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_512
timestamp 1666464484
transform 1 0 58688 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_522
timestamp 1666464484
transform 1 0 59808 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_532
timestamp 1666464484
transform 1 0 60928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_542
timestamp 1666464484
transform 1 0 62048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_544
timestamp 1666464484
transform 1 0 62272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_551
timestamp 1666464484
transform 1 0 63056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_559
timestamp 1666464484
transform 1 0 63952 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1666464484
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_570
timestamp 1666464484
transform 1 0 65184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_575
timestamp 1666464484
transform 1 0 65744 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_585
timestamp 1666464484
transform 1 0 66864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_596
timestamp 1666464484
transform 1 0 68096 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_609
timestamp 1666464484
transform 1 0 69552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_623
timestamp 1666464484
transform 1 0 71120 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1666464484
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_641
timestamp 1666464484
transform 1 0 73136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_656
timestamp 1666464484
transform 1 0 74816 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_664
timestamp 1666464484
transform 1 0 75712 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_678
timestamp 1666464484
transform 1 0 77280 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_688
timestamp 1666464484
transform 1 0 78400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_696
timestamp 1666464484
transform 1 0 79296 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_702
timestamp 1666464484
transform 1 0 79968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_709
timestamp 1666464484
transform 1 0 80752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_712
timestamp 1666464484
transform 1 0 81088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_718
timestamp 1666464484
transform 1 0 81760 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_729
timestamp 1666464484
transform 1 0 82992 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_731
timestamp 1666464484
transform 1 0 83216 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_769
timestamp 1666464484
transform 1 0 87472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_777
timestamp 1666464484
transform 1 0 88368 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_783
timestamp 1666464484
transform 1 0 89040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_786
timestamp 1666464484
transform 1 0 89376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_802
timestamp 1666464484
transform 1 0 91168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_810
timestamp 1666464484
transform 1 0 92064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_817
timestamp 1666464484
transform 1 0 92848 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_821
timestamp 1666464484
transform 1 0 93296 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_825
timestamp 1666464484
transform 1 0 93744 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_829
timestamp 1666464484
transform 1 0 94192 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_831
timestamp 1666464484
transform 1 0 94416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_838
timestamp 1666464484
transform 1 0 95200 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_851
timestamp 1666464484
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_854
timestamp 1666464484
transform 1 0 96992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_868
timestamp 1666464484
transform 1 0 98560 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_876
timestamp 1666464484
transform 1 0 99456 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_884
timestamp 1666464484
transform 1 0 100352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_888
timestamp 1666464484
transform 1 0 100800 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_890
timestamp 1666464484
transform 1 0 101024 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_901
timestamp 1666464484
transform 1 0 102256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_905
timestamp 1666464484
transform 1 0 102704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_911
timestamp 1666464484
transform 1 0 103376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_915
timestamp 1666464484
transform 1 0 103824 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_922
timestamp 1666464484
transform 1 0 104608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_925
timestamp 1666464484
transform 1 0 104944 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_939
timestamp 1666464484
transform 1 0 106512 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_949
timestamp 1666464484
transform 1 0 107632 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_957
timestamp 1666464484
transform 1 0 108528 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_992
timestamp 1666464484
transform 1 0 112448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_996
timestamp 1666464484
transform 1 0 112896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1007
timestamp 1666464484
transform 1 0 114128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1011
timestamp 1666464484
transform 1 0 114576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1015
timestamp 1666464484
transform 1 0 115024 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1022
timestamp 1666464484
transform 1 0 115808 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1026
timestamp 1666464484
transform 1 0 116256 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1030
timestamp 1666464484
transform 1 0 116704 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1034
timestamp 1666464484
transform 1 0 117152 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1036
timestamp 1666464484
transform 1 0 117376 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1041
timestamp 1666464484
transform 1 0 117936 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1051
timestamp 1666464484
transform 1 0 119056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1061
timestamp 1666464484
transform 1 0 120176 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1067
timestamp 1666464484
transform 1 0 120848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1074
timestamp 1666464484
transform 1 0 121632 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1082
timestamp 1666464484
transform 1 0 122528 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1090
timestamp 1666464484
transform 1 0 123424 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1098
timestamp 1666464484
transform 1 0 124320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1106
timestamp 1666464484
transform 1 0 125216 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1110
timestamp 1666464484
transform 1 0 125664 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1114
timestamp 1666464484
transform 1 0 126112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1118
timestamp 1666464484
transform 1 0 126560 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1122
timestamp 1666464484
transform 1 0 127008 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1126
timestamp 1666464484
transform 1 0 127456 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1128
timestamp 1666464484
transform 1 0 127680 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1135
timestamp 1666464484
transform 1 0 128464 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1138
timestamp 1666464484
transform 1 0 128800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1145
timestamp 1666464484
transform 1 0 129584 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1153
timestamp 1666464484
transform 1 0 130480 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1161
timestamp 1666464484
transform 1 0 131376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1167
timestamp 1666464484
transform 1 0 132048 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1177
timestamp 1666464484
transform 1 0 133168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1179
timestamp 1666464484
transform 1 0 133392 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1186
timestamp 1666464484
transform 1 0 134176 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1194
timestamp 1666464484
transform 1 0 135072 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1202
timestamp 1666464484
transform 1 0 135968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1206
timestamp 1666464484
transform 1 0 136416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1209
timestamp 1666464484
transform 1 0 136752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1216
timestamp 1666464484
transform 1 0 137536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1220
timestamp 1666464484
transform 1 0 137984 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1226
timestamp 1666464484
transform 1 0 138656 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1230
timestamp 1666464484
transform 1 0 139104 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1234
timestamp 1666464484
transform 1 0 139552 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1241
timestamp 1666464484
transform 1 0 140336 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1249
timestamp 1666464484
transform 1 0 141232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1251
timestamp 1666464484
transform 1 0 141456 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1256
timestamp 1666464484
transform 1 0 142016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1264
timestamp 1666464484
transform 1 0 142912 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1266
timestamp 1666464484
transform 1 0 143136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1271
timestamp 1666464484
transform 1 0 143696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1275
timestamp 1666464484
transform 1 0 144144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1277
timestamp 1666464484
transform 1 0 144368 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1280
timestamp 1666464484
transform 1 0 144704 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1290
timestamp 1666464484
transform 1 0 145824 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1294
timestamp 1666464484
transform 1 0 146272 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1296
timestamp 1666464484
transform 1 0 146496 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1301
timestamp 1666464484
transform 1 0 147056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1305
timestamp 1666464484
transform 1 0 147504 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1309
timestamp 1666464484
transform 1 0 147952 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1313
timestamp 1666464484
transform 1 0 148400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1317
timestamp 1666464484
transform 1 0 148848 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1321
timestamp 1666464484
transform 1 0 149296 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1325
timestamp 1666464484
transform 1 0 149744 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1329
timestamp 1666464484
transform 1 0 150192 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1345
timestamp 1666464484
transform 1 0 151984 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1351 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 152656 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1415
timestamp 1666464484
transform 1 0 159824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1419
timestamp 1666464484
transform 1 0 160272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1422
timestamp 1666464484
transform 1 0 160608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1486
timestamp 1666464484
transform 1 0 167776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1490
timestamp 1666464484
transform 1 0 168224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_1493
timestamp 1666464484
transform 1 0 168560 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1557
timestamp 1666464484
transform 1 0 175728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1561
timestamp 1666464484
transform 1 0 176176 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1564
timestamp 1666464484
transform 1 0 176512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1580
timestamp 1666464484
transform 1 0 178304 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1666464484
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1666464484
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1666464484
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1666464484
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_108
timestamp 1666464484
transform 1 0 13440 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_112
timestamp 1666464484
transform 1 0 13888 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_115
timestamp 1666464484
transform 1 0 14224 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_123
timestamp 1666464484
transform 1 0 15120 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_127
timestamp 1666464484
transform 1 0 15568 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_131
timestamp 1666464484
transform 1 0 16016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_135
timestamp 1666464484
transform 1 0 16464 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_137
timestamp 1666464484
transform 1 0 16688 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_140
timestamp 1666464484
transform 1 0 17024 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_144
timestamp 1666464484
transform 1 0 17472 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_148
timestamp 1666464484
transform 1 0 17920 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_152
timestamp 1666464484
transform 1 0 18368 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_159
timestamp 1666464484
transform 1 0 19152 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1666464484
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1666464484
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_182
timestamp 1666464484
transform 1 0 21728 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_184
timestamp 1666464484
transform 1 0 21952 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_187
timestamp 1666464484
transform 1 0 22288 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_197
timestamp 1666464484
transform 1 0 23408 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_207
timestamp 1666464484
transform 1 0 24528 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_211
timestamp 1666464484
transform 1 0 24976 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_215
timestamp 1666464484
transform 1 0 25424 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_223
timestamp 1666464484
transform 1 0 26320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_229
timestamp 1666464484
transform 1 0 26992 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_246
timestamp 1666464484
transform 1 0 28896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1666464484
transform 1 0 29344 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_257
timestamp 1666464484
transform 1 0 30128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_267
timestamp 1666464484
transform 1 0 31248 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_271
timestamp 1666464484
transform 1 0 31696 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_302
timestamp 1666464484
transform 1 0 35168 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_314
timestamp 1666464484
transform 1 0 36512 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1666464484
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_321
timestamp 1666464484
transform 1 0 37296 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_330
timestamp 1666464484
transform 1 0 38304 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_332
timestamp 1666464484
transform 1 0 38528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_339
timestamp 1666464484
transform 1 0 39312 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_347
timestamp 1666464484
transform 1 0 40208 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_355
timestamp 1666464484
transform 1 0 41104 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_363
timestamp 1666464484
transform 1 0 42000 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_376
timestamp 1666464484
transform 1 0 43456 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_378
timestamp 1666464484
transform 1 0 43680 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_381
timestamp 1666464484
transform 1 0 44016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1666464484
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1666464484
transform 1 0 45248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_408
timestamp 1666464484
transform 1 0 47040 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_412
timestamp 1666464484
transform 1 0 47488 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_419
timestamp 1666464484
transform 1 0 48272 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_427
timestamp 1666464484
transform 1 0 49168 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_444
timestamp 1666464484
transform 1 0 51072 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1666464484
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_463
timestamp 1666464484
transform 1 0 53200 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_493
timestamp 1666464484
transform 1 0 56560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_497
timestamp 1666464484
transform 1 0 57008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_500
timestamp 1666464484
transform 1 0 57344 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_508
timestamp 1666464484
transform 1 0 58240 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_512
timestamp 1666464484
transform 1 0 58688 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_515
timestamp 1666464484
transform 1 0 59024 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_523
timestamp 1666464484
transform 1 0 59920 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_534
timestamp 1666464484
transform 1 0 61152 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_540
timestamp 1666464484
transform 1 0 61824 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_571
timestamp 1666464484
transform 1 0 65296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_575
timestamp 1666464484
transform 1 0 65744 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_589
timestamp 1666464484
transform 1 0 67312 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_598
timestamp 1666464484
transform 1 0 68320 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1666464484
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_605
timestamp 1666464484
transform 1 0 69104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_656
timestamp 1666464484
transform 1 0 74816 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_664
timestamp 1666464484
transform 1 0 75712 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_666
timestamp 1666464484
transform 1 0 75936 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1666464484
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_676
timestamp 1666464484
transform 1 0 77056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_685
timestamp 1666464484
transform 1 0 78064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_693
timestamp 1666464484
transform 1 0 78960 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_697
timestamp 1666464484
transform 1 0 79408 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_703
timestamp 1666464484
transform 1 0 80080 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_717
timestamp 1666464484
transform 1 0 81648 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_719
timestamp 1666464484
transform 1 0 81872 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_725
timestamp 1666464484
transform 1 0 82544 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_735
timestamp 1666464484
transform 1 0 83664 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_737
timestamp 1666464484
transform 1 0 83888 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1666464484
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_747
timestamp 1666464484
transform 1 0 85008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_757
timestamp 1666464484
transform 1 0 86128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_765
timestamp 1666464484
transform 1 0 87024 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_769
timestamp 1666464484
transform 1 0 87472 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_773
timestamp 1666464484
transform 1 0 87920 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_779
timestamp 1666464484
transform 1 0 88592 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_783
timestamp 1666464484
transform 1 0 89040 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_786
timestamp 1666464484
transform 1 0 89376 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_790
timestamp 1666464484
transform 1 0 89824 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_794
timestamp 1666464484
transform 1 0 90272 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_798
timestamp 1666464484
transform 1 0 90720 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_802
timestamp 1666464484
transform 1 0 91168 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_806
timestamp 1666464484
transform 1 0 91616 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_810
timestamp 1666464484
transform 1 0 92064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_814
timestamp 1666464484
transform 1 0 92512 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_818
timestamp 1666464484
transform 1 0 92960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_821
timestamp 1666464484
transform 1 0 93296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_827
timestamp 1666464484
transform 1 0 93968 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_829
timestamp 1666464484
transform 1 0 94192 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_832
timestamp 1666464484
transform 1 0 94528 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_836
timestamp 1666464484
transform 1 0 94976 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_839
timestamp 1666464484
transform 1 0 95312 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_849
timestamp 1666464484
transform 1 0 96432 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_853
timestamp 1666464484
transform 1 0 96880 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_862
timestamp 1666464484
transform 1 0 97888 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_870
timestamp 1666464484
transform 1 0 98784 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_874
timestamp 1666464484
transform 1 0 99232 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_878
timestamp 1666464484
transform 1 0 99680 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_882
timestamp 1666464484
transform 1 0 100128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_886
timestamp 1666464484
transform 1 0 100576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_889
timestamp 1666464484
transform 1 0 100912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_892
timestamp 1666464484
transform 1 0 101248 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_896
timestamp 1666464484
transform 1 0 101696 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_910
timestamp 1666464484
transform 1 0 103264 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_914
timestamp 1666464484
transform 1 0 103712 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_923
timestamp 1666464484
transform 1 0 104720 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_957
timestamp 1666464484
transform 1 0 108528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_960
timestamp 1666464484
transform 1 0 108864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_967
timestamp 1666464484
transform 1 0 109648 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_977
timestamp 1666464484
transform 1 0 110768 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_983
timestamp 1666464484
transform 1 0 111440 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_987
timestamp 1666464484
transform 1 0 111888 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_991
timestamp 1666464484
transform 1 0 112336 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_995
timestamp 1666464484
transform 1 0 112784 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_999
timestamp 1666464484
transform 1 0 113232 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1003
timestamp 1666464484
transform 1 0 113680 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1007
timestamp 1666464484
transform 1 0 114128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1011
timestamp 1666464484
transform 1 0 114576 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1015
timestamp 1666464484
transform 1 0 115024 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1017
timestamp 1666464484
transform 1 0 115248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1028
timestamp 1666464484
transform 1 0 116480 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1031
timestamp 1666464484
transform 1 0 116816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1034
timestamp 1666464484
transform 1 0 117152 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1038
timestamp 1666464484
transform 1 0 117600 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1042
timestamp 1666464484
transform 1 0 118048 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1046
timestamp 1666464484
transform 1 0 118496 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1055
timestamp 1666464484
transform 1 0 119504 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1071
timestamp 1666464484
transform 1 0 121296 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1075
timestamp 1666464484
transform 1 0 121744 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1079
timestamp 1666464484
transform 1 0 122192 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1083
timestamp 1666464484
transform 1 0 122640 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1087
timestamp 1666464484
transform 1 0 123088 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1091
timestamp 1666464484
transform 1 0 123536 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1095
timestamp 1666464484
transform 1 0 123984 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1099
timestamp 1666464484
transform 1 0 124432 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1102
timestamp 1666464484
transform 1 0 124768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1105
timestamp 1666464484
transform 1 0 125104 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1109
timestamp 1666464484
transform 1 0 125552 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1113
timestamp 1666464484
transform 1 0 126000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1119
timestamp 1666464484
transform 1 0 126672 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1123
timestamp 1666464484
transform 1 0 127120 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1127
timestamp 1666464484
transform 1 0 127568 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1133
timestamp 1666464484
transform 1 0 128240 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1137
timestamp 1666464484
transform 1 0 128688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1141
timestamp 1666464484
transform 1 0 129136 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1151
timestamp 1666464484
transform 1 0 130256 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1159
timestamp 1666464484
transform 1 0 131152 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1161
timestamp 1666464484
transform 1 0 131376 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1166
timestamp 1666464484
transform 1 0 131936 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1170
timestamp 1666464484
transform 1 0 132384 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1173
timestamp 1666464484
transform 1 0 132720 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1181
timestamp 1666464484
transform 1 0 133616 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1185
timestamp 1666464484
transform 1 0 134064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1189
timestamp 1666464484
transform 1 0 134512 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1191
timestamp 1666464484
transform 1 0 134736 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1196
timestamp 1666464484
transform 1 0 135296 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1198
timestamp 1666464484
transform 1 0 135520 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1205
timestamp 1666464484
transform 1 0 136304 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1211
timestamp 1666464484
transform 1 0 136976 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1215
timestamp 1666464484
transform 1 0 137424 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1219
timestamp 1666464484
transform 1 0 137872 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1223
timestamp 1666464484
transform 1 0 138320 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1227
timestamp 1666464484
transform 1 0 138768 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1231
timestamp 1666464484
transform 1 0 139216 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1235
timestamp 1666464484
transform 1 0 139664 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1239
timestamp 1666464484
transform 1 0 140112 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1241
timestamp 1666464484
transform 1 0 140336 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1244
timestamp 1666464484
transform 1 0 140672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1247
timestamp 1666464484
transform 1 0 141008 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1251
timestamp 1666464484
transform 1 0 141456 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1255
timestamp 1666464484
transform 1 0 141904 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1259
timestamp 1666464484
transform 1 0 142352 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1263
timestamp 1666464484
transform 1 0 142800 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1267
timestamp 1666464484
transform 1 0 143248 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1271
timestamp 1666464484
transform 1 0 143696 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1275
timestamp 1666464484
transform 1 0 144144 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1277
timestamp 1666464484
transform 1 0 144368 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1280
timestamp 1666464484
transform 1 0 144704 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1286
timestamp 1666464484
transform 1 0 145376 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1288
timestamp 1666464484
transform 1 0 145600 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1291
timestamp 1666464484
transform 1 0 145936 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1295
timestamp 1666464484
transform 1 0 146384 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1299
timestamp 1666464484
transform 1 0 146832 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1303
timestamp 1666464484
transform 1 0 147280 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1307
timestamp 1666464484
transform 1 0 147728 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1311
timestamp 1666464484
transform 1 0 148176 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1315
timestamp 1666464484
transform 1 0 148624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1318
timestamp 1666464484
transform 1 0 148960 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1382
timestamp 1666464484
transform 1 0 156128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1386
timestamp 1666464484
transform 1 0 156576 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1450
timestamp 1666464484
transform 1 0 163744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1454
timestamp 1666464484
transform 1 0 164192 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_1457
timestamp 1666464484
transform 1 0 164528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1521
timestamp 1666464484
transform 1 0 171696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1525
timestamp 1666464484
transform 1 0 172144 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1528
timestamp 1666464484
transform 1 0 172480 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1560
timestamp 1666464484
transform 1 0 176064 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1576
timestamp 1666464484
transform 1 0 177856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1580
timestamp 1666464484
transform 1 0 178304 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1666464484
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1666464484
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_73
timestamp 1666464484
transform 1 0 9520 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_105
timestamp 1666464484
transform 1 0 13104 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_113
timestamp 1666464484
transform 1 0 14000 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_117
timestamp 1666464484
transform 1 0 14448 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_119
timestamp 1666464484
transform 1 0 14672 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_122
timestamp 1666464484
transform 1 0 15008 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_130
timestamp 1666464484
transform 1 0 15904 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_132
timestamp 1666464484
transform 1 0 16128 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_135
timestamp 1666464484
transform 1 0 16464 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_139
timestamp 1666464484
transform 1 0 16912 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1666464484
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_144
timestamp 1666464484
transform 1 0 17472 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_148
timestamp 1666464484
transform 1 0 17920 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_178
timestamp 1666464484
transform 1 0 21280 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_182
timestamp 1666464484
transform 1 0 21728 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_186
timestamp 1666464484
transform 1 0 22176 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_190
timestamp 1666464484
transform 1 0 22624 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_194
timestamp 1666464484
transform 1 0 23072 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_198
timestamp 1666464484
transform 1 0 23520 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_202
timestamp 1666464484
transform 1 0 23968 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1666464484
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_210
timestamp 1666464484
transform 1 0 24864 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1666464484
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1666464484
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_245
timestamp 1666464484
transform 1 0 28784 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_249
timestamp 1666464484
transform 1 0 29232 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_253
timestamp 1666464484
transform 1 0 29680 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_257
timestamp 1666464484
transform 1 0 30128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_259
timestamp 1666464484
transform 1 0 30352 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_262
timestamp 1666464484
transform 1 0 30688 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_266
timestamp 1666464484
transform 1 0 31136 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_270
timestamp 1666464484
transform 1 0 31584 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_278
timestamp 1666464484
transform 1 0 32480 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_280
timestamp 1666464484
transform 1 0 32704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1666464484
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_286
timestamp 1666464484
transform 1 0 33376 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_289
timestamp 1666464484
transform 1 0 33712 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_299
timestamp 1666464484
transform 1 0 34832 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_301
timestamp 1666464484
transform 1 0 35056 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_304
timestamp 1666464484
transform 1 0 35392 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_312
timestamp 1666464484
transform 1 0 36288 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_316
timestamp 1666464484
transform 1 0 36736 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_320
timestamp 1666464484
transform 1 0 37184 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_328
timestamp 1666464484
transform 1 0 38080 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_332
timestamp 1666464484
transform 1 0 38528 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_335
timestamp 1666464484
transform 1 0 38864 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_343
timestamp 1666464484
transform 1 0 39760 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_347
timestamp 1666464484
transform 1 0 40208 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_350
timestamp 1666464484
transform 1 0 40544 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1666464484
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_357
timestamp 1666464484
transform 1 0 41328 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_360
timestamp 1666464484
transform 1 0 41664 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_364
timestamp 1666464484
transform 1 0 42112 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_372
timestamp 1666464484
transform 1 0 43008 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_403
timestamp 1666464484
transform 1 0 46480 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_405
timestamp 1666464484
transform 1 0 46704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_412
timestamp 1666464484
transform 1 0 47488 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_422
timestamp 1666464484
transform 1 0 48608 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1666464484
transform 1 0 49280 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_479
timestamp 1666464484
transform 1 0 54992 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_487
timestamp 1666464484
transform 1 0 55888 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_489
timestamp 1666464484
transform 1 0 56112 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1666464484
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_499
timestamp 1666464484
transform 1 0 57232 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_532
timestamp 1666464484
transform 1 0 60928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_534
timestamp 1666464484
transform 1 0 61152 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_537
timestamp 1666464484
transform 1 0 61488 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_541
timestamp 1666464484
transform 1 0 61936 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_551
timestamp 1666464484
transform 1 0 63056 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_561
timestamp 1666464484
transform 1 0 64176 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1666464484
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_570
timestamp 1666464484
transform 1 0 65184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_621
timestamp 1666464484
transform 1 0 70896 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_623
timestamp 1666464484
transform 1 0 71120 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_637
timestamp 1666464484
transform 1 0 72688 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_641
timestamp 1666464484
transform 1 0 73136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_648
timestamp 1666464484
transform 1 0 73920 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_656
timestamp 1666464484
transform 1 0 74816 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_658
timestamp 1666464484
transform 1 0 75040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_664
timestamp 1666464484
transform 1 0 75712 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_668
timestamp 1666464484
transform 1 0 76160 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_706
timestamp 1666464484
transform 1 0 80416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_712
timestamp 1666464484
transform 1 0 81088 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_714
timestamp 1666464484
transform 1 0 81312 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_720
timestamp 1666464484
transform 1 0 81984 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_754
timestamp 1666464484
transform 1 0 85792 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_756
timestamp 1666464484
transform 1 0 86016 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_769
timestamp 1666464484
transform 1 0 87472 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_773
timestamp 1666464484
transform 1 0 87920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_777
timestamp 1666464484
transform 1 0 88368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1666464484
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_783
timestamp 1666464484
transform 1 0 89040 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_797
timestamp 1666464484
transform 1 0 90608 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_801
timestamp 1666464484
transform 1 0 91056 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_805
timestamp 1666464484
transform 1 0 91504 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_808
timestamp 1666464484
transform 1 0 91840 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_812
timestamp 1666464484
transform 1 0 92288 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_814
timestamp 1666464484
transform 1 0 92512 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_817
timestamp 1666464484
transform 1 0 92848 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_821
timestamp 1666464484
transform 1 0 93296 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_825
timestamp 1666464484
transform 1 0 93744 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_829
timestamp 1666464484
transform 1 0 94192 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_833
timestamp 1666464484
transform 1 0 94640 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_844
timestamp 1666464484
transform 1 0 95872 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_848
timestamp 1666464484
transform 1 0 96320 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_854
timestamp 1666464484
transform 1 0 96992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_859
timestamp 1666464484
transform 1 0 97552 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_863
timestamp 1666464484
transform 1 0 98000 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_867
timestamp 1666464484
transform 1 0 98448 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_871
timestamp 1666464484
transform 1 0 98896 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_875
timestamp 1666464484
transform 1 0 99344 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_879
timestamp 1666464484
transform 1 0 99792 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_883
timestamp 1666464484
transform 1 0 100240 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_887
timestamp 1666464484
transform 1 0 100688 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_891
timestamp 1666464484
transform 1 0 101136 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_899
timestamp 1666464484
transform 1 0 102032 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_907
timestamp 1666464484
transform 1 0 102928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_915
timestamp 1666464484
transform 1 0 103824 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_921
timestamp 1666464484
transform 1 0 104496 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_925
timestamp 1666464484
transform 1 0 104944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_928
timestamp 1666464484
transform 1 0 105280 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_932
timestamp 1666464484
transform 1 0 105728 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_936
timestamp 1666464484
transform 1 0 106176 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_940
timestamp 1666464484
transform 1 0 106624 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_944
timestamp 1666464484
transform 1 0 107072 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_948
timestamp 1666464484
transform 1 0 107520 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_955
timestamp 1666464484
transform 1 0 108304 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_959
timestamp 1666464484
transform 1 0 108752 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_963
timestamp 1666464484
transform 1 0 109200 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_967
timestamp 1666464484
transform 1 0 109648 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_971
timestamp 1666464484
transform 1 0 110096 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_975
timestamp 1666464484
transform 1 0 110544 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_979
timestamp 1666464484
transform 1 0 110992 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_983
timestamp 1666464484
transform 1 0 111440 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_993
timestamp 1666464484
transform 1 0 112560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_996
timestamp 1666464484
transform 1 0 112896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1003
timestamp 1666464484
transform 1 0 113680 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1007
timestamp 1666464484
transform 1 0 114128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1011
timestamp 1666464484
transform 1 0 114576 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1015
timestamp 1666464484
transform 1 0 115024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1025
timestamp 1666464484
transform 1 0 116144 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1029
timestamp 1666464484
transform 1 0 116592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1033
timestamp 1666464484
transform 1 0 117040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1040
timestamp 1666464484
transform 1 0 117824 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1050
timestamp 1666464484
transform 1 0 118944 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1064
timestamp 1666464484
transform 1 0 120512 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1067
timestamp 1666464484
transform 1 0 120848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1070
timestamp 1666464484
transform 1 0 121184 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1074
timestamp 1666464484
transform 1 0 121632 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1078
timestamp 1666464484
transform 1 0 122080 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1082
timestamp 1666464484
transform 1 0 122528 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1086
timestamp 1666464484
transform 1 0 122976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1090
timestamp 1666464484
transform 1 0 123424 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1094
timestamp 1666464484
transform 1 0 123872 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1098
timestamp 1666464484
transform 1 0 124320 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1102
timestamp 1666464484
transform 1 0 124768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1106
timestamp 1666464484
transform 1 0 125216 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1110
timestamp 1666464484
transform 1 0 125664 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1112
timestamp 1666464484
transform 1 0 125888 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1115
timestamp 1666464484
transform 1 0 126224 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1119
timestamp 1666464484
transform 1 0 126672 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1127
timestamp 1666464484
transform 1 0 127568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1131
timestamp 1666464484
transform 1 0 128016 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1135
timestamp 1666464484
transform 1 0 128464 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1138
timestamp 1666464484
transform 1 0 128800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1141
timestamp 1666464484
transform 1 0 129136 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1145
timestamp 1666464484
transform 1 0 129584 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1149
timestamp 1666464484
transform 1 0 130032 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1153
timestamp 1666464484
transform 1 0 130480 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1157
timestamp 1666464484
transform 1 0 130928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1163
timestamp 1666464484
transform 1 0 131600 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1167
timestamp 1666464484
transform 1 0 132048 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1171
timestamp 1666464484
transform 1 0 132496 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1175
timestamp 1666464484
transform 1 0 132944 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1179
timestamp 1666464484
transform 1 0 133392 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1183
timestamp 1666464484
transform 1 0 133840 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1186
timestamp 1666464484
transform 1 0 134176 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1190
timestamp 1666464484
transform 1 0 134624 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1196
timestamp 1666464484
transform 1 0 135296 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1200
timestamp 1666464484
transform 1 0 135744 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1204
timestamp 1666464484
transform 1 0 136192 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1206
timestamp 1666464484
transform 1 0 136416 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1209
timestamp 1666464484
transform 1 0 136752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1212
timestamp 1666464484
transform 1 0 137088 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1216
timestamp 1666464484
transform 1 0 137536 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1220
timestamp 1666464484
transform 1 0 137984 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1224
timestamp 1666464484
transform 1 0 138432 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1228
timestamp 1666464484
transform 1 0 138880 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1232
timestamp 1666464484
transform 1 0 139328 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1236
timestamp 1666464484
transform 1 0 139776 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1239
timestamp 1666464484
transform 1 0 140112 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1243
timestamp 1666464484
transform 1 0 140560 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1247
timestamp 1666464484
transform 1 0 141008 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1253
timestamp 1666464484
transform 1 0 141680 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1257
timestamp 1666464484
transform 1 0 142128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1263
timestamp 1666464484
transform 1 0 142800 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1267
timestamp 1666464484
transform 1 0 143248 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1271
timestamp 1666464484
transform 1 0 143696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1275
timestamp 1666464484
transform 1 0 144144 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1277
timestamp 1666464484
transform 1 0 144368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1280
timestamp 1666464484
transform 1 0 144704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1283
timestamp 1666464484
transform 1 0 145040 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1287
timestamp 1666464484
transform 1 0 145488 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1319
timestamp 1666464484
transform 1 0 149072 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1335
timestamp 1666464484
transform 1 0 150864 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1343
timestamp 1666464484
transform 1 0 151760 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1347
timestamp 1666464484
transform 1 0 152208 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1351
timestamp 1666464484
transform 1 0 152656 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1415
timestamp 1666464484
transform 1 0 159824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1419
timestamp 1666464484
transform 1 0 160272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1422
timestamp 1666464484
transform 1 0 160608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1486
timestamp 1666464484
transform 1 0 167776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1490
timestamp 1666464484
transform 1 0 168224 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1493
timestamp 1666464484
transform 1 0 168560 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1557
timestamp 1666464484
transform 1 0 175728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1561
timestamp 1666464484
transform 1 0 176176 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1564
timestamp 1666464484
transform 1 0 176512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1580
timestamp 1666464484
transform 1 0 178304 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1666464484
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1666464484
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1666464484
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1666464484
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1666464484
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_108
timestamp 1666464484
transform 1 0 13440 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_140
timestamp 1666464484
transform 1 0 17024 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_156
timestamp 1666464484
transform 1 0 18816 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_158
timestamp 1666464484
transform 1 0 19040 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_165
timestamp 1666464484
transform 1 0 19824 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_173
timestamp 1666464484
transform 1 0 20720 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_179
timestamp 1666464484
transform 1 0 21392 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_211
timestamp 1666464484
transform 1 0 24976 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_219
timestamp 1666464484
transform 1 0 25872 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_223
timestamp 1666464484
transform 1 0 26320 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_225
timestamp 1666464484
transform 1 0 26544 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_232
timestamp 1666464484
transform 1 0 27328 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_238
timestamp 1666464484
transform 1 0 28000 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_242
timestamp 1666464484
transform 1 0 28448 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_244
timestamp 1666464484
transform 1 0 28672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1666464484
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_250
timestamp 1666464484
transform 1 0 29344 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_253
timestamp 1666464484
transform 1 0 29680 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_290
timestamp 1666464484
transform 1 0 33824 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_307
timestamp 1666464484
transform 1 0 35728 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_311
timestamp 1666464484
transform 1 0 36176 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_314
timestamp 1666464484
transform 1 0 36512 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1666464484
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_321
timestamp 1666464484
transform 1 0 37296 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_323
timestamp 1666464484
transform 1 0 37520 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_339
timestamp 1666464484
transform 1 0 39312 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_356
timestamp 1666464484
transform 1 0 41216 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_362
timestamp 1666464484
transform 1 0 41888 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_366
timestamp 1666464484
transform 1 0 42336 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_370
timestamp 1666464484
transform 1 0 42784 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_374
timestamp 1666464484
transform 1 0 43232 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_382
timestamp 1666464484
transform 1 0 44128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_386
timestamp 1666464484
transform 1 0 44576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1666464484
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_392
timestamp 1666464484
transform 1 0 45248 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_399
timestamp 1666464484
transform 1 0 46032 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_407
timestamp 1666464484
transform 1 0 46928 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_415
timestamp 1666464484
transform 1 0 47824 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_446
timestamp 1666464484
transform 1 0 51296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_458
timestamp 1666464484
transform 1 0 52640 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1666464484
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_463
timestamp 1666464484
transform 1 0 53200 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_472
timestamp 1666464484
transform 1 0 54208 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_484
timestamp 1666464484
transform 1 0 55552 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_492
timestamp 1666464484
transform 1 0 56448 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_498
timestamp 1666464484
transform 1 0 57120 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_506
timestamp 1666464484
transform 1 0 58016 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_508
timestamp 1666464484
transform 1 0 58240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_511
timestamp 1666464484
transform 1 0 58576 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_515
timestamp 1666464484
transform 1 0 59024 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_519
timestamp 1666464484
transform 1 0 59472 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_523
timestamp 1666464484
transform 1 0 59920 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_527
timestamp 1666464484
transform 1 0 60368 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_534
timestamp 1666464484
transform 1 0 61152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_585
timestamp 1666464484
transform 1 0 66864 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_587
timestamp 1666464484
transform 1 0 67088 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_594
timestamp 1666464484
transform 1 0 67872 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1666464484
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_605
timestamp 1666464484
transform 1 0 69104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_656
timestamp 1666464484
transform 1 0 74816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_665
timestamp 1666464484
transform 1 0 75824 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1666464484
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_676
timestamp 1666464484
transform 1 0 77056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_683
timestamp 1666464484
transform 1 0 77840 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_691
timestamp 1666464484
transform 1 0 78736 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_698
timestamp 1666464484
transform 1 0 79520 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_706
timestamp 1666464484
transform 1 0 80416 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_716
timestamp 1666464484
transform 1 0 81536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_720
timestamp 1666464484
transform 1 0 81984 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_733
timestamp 1666464484
transform 1 0 83440 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_737
timestamp 1666464484
transform 1 0 83888 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1666464484
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_747
timestamp 1666464484
transform 1 0 85008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_756
timestamp 1666464484
transform 1 0 86016 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_760
timestamp 1666464484
transform 1 0 86464 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_764
timestamp 1666464484
transform 1 0 86912 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_774
timestamp 1666464484
transform 1 0 88032 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_782
timestamp 1666464484
transform 1 0 88928 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_788
timestamp 1666464484
transform 1 0 89600 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_803
timestamp 1666464484
transform 1 0 91280 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_811
timestamp 1666464484
transform 1 0 92176 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1666464484
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_818
timestamp 1666464484
transform 1 0 92960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_821
timestamp 1666464484
transform 1 0 93296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_827
timestamp 1666464484
transform 1 0 93968 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_831
timestamp 1666464484
transform 1 0 94416 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_844
timestamp 1666464484
transform 1 0 95872 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_854
timestamp 1666464484
transform 1 0 96992 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_858
timestamp 1666464484
transform 1 0 97440 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_871
timestamp 1666464484
transform 1 0 98896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_880
timestamp 1666464484
transform 1 0 99904 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_884
timestamp 1666464484
transform 1 0 100352 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1666464484
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_889
timestamp 1666464484
transform 1 0 100912 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_891
timestamp 1666464484
transform 1 0 101136 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_900
timestamp 1666464484
transform 1 0 102144 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_904
timestamp 1666464484
transform 1 0 102592 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_908
timestamp 1666464484
transform 1 0 103040 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_918
timestamp 1666464484
transform 1 0 104160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_922
timestamp 1666464484
transform 1 0 104608 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_930
timestamp 1666464484
transform 1 0 105504 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_934
timestamp 1666464484
transform 1 0 105952 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_938
timestamp 1666464484
transform 1 0 106400 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_942
timestamp 1666464484
transform 1 0 106848 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_946
timestamp 1666464484
transform 1 0 107296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_950
timestamp 1666464484
transform 1 0 107744 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_957
timestamp 1666464484
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_960
timestamp 1666464484
transform 1 0 108864 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_993
timestamp 1666464484
transform 1 0 112560 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_997
timestamp 1666464484
transform 1 0 113008 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1001
timestamp 1666464484
transform 1 0 113456 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1005
timestamp 1666464484
transform 1 0 113904 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1009
timestamp 1666464484
transform 1 0 114352 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1011
timestamp 1666464484
transform 1 0 114576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1018
timestamp 1666464484
transform 1 0 115360 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1026
timestamp 1666464484
transform 1 0 116256 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1028
timestamp 1666464484
transform 1 0 116480 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1031
timestamp 1666464484
transform 1 0 116816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1034
timestamp 1666464484
transform 1 0 117152 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1038
timestamp 1666464484
transform 1 0 117600 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1042
timestamp 1666464484
transform 1 0 118048 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1046
timestamp 1666464484
transform 1 0 118496 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1050
timestamp 1666464484
transform 1 0 118944 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1052
timestamp 1666464484
transform 1 0 119168 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1063
timestamp 1666464484
transform 1 0 120400 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1067
timestamp 1666464484
transform 1 0 120848 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1071
timestamp 1666464484
transform 1 0 121296 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1075
timestamp 1666464484
transform 1 0 121744 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1079
timestamp 1666464484
transform 1 0 122192 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1083
timestamp 1666464484
transform 1 0 122640 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1087
timestamp 1666464484
transform 1 0 123088 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1091
timestamp 1666464484
transform 1 0 123536 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1095
timestamp 1666464484
transform 1 0 123984 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1099
timestamp 1666464484
transform 1 0 124432 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1102
timestamp 1666464484
transform 1 0 124768 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1134
timestamp 1666464484
transform 1 0 128352 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1136
timestamp 1666464484
transform 1 0 128576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1139
timestamp 1666464484
transform 1 0 128912 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1147
timestamp 1666464484
transform 1 0 129808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1151
timestamp 1666464484
transform 1 0 130256 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1155
timestamp 1666464484
transform 1 0 130704 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1159
timestamp 1666464484
transform 1 0 131152 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1163
timestamp 1666464484
transform 1 0 131600 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1167
timestamp 1666464484
transform 1 0 132048 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1173
timestamp 1666464484
transform 1 0 132720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1176
timestamp 1666464484
transform 1 0 133056 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1182
timestamp 1666464484
transform 1 0 133728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1190
timestamp 1666464484
transform 1 0 134624 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1192
timestamp 1666464484
transform 1 0 134848 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1195
timestamp 1666464484
transform 1 0 135184 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1199
timestamp 1666464484
transform 1 0 135632 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1209
timestamp 1666464484
transform 1 0 136752 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1213
timestamp 1666464484
transform 1 0 137200 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1217
timestamp 1666464484
transform 1 0 137648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1225
timestamp 1666464484
transform 1 0 138544 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1228
timestamp 1666464484
transform 1 0 138880 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1232
timestamp 1666464484
transform 1 0 139328 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1236
timestamp 1666464484
transform 1 0 139776 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1240
timestamp 1666464484
transform 1 0 140224 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1244
timestamp 1666464484
transform 1 0 140672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1247
timestamp 1666464484
transform 1 0 141008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1311
timestamp 1666464484
transform 1 0 148176 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1315
timestamp 1666464484
transform 1 0 148624 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1379
timestamp 1666464484
transform 1 0 155792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1383
timestamp 1666464484
transform 1 0 156240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1386
timestamp 1666464484
transform 1 0 156576 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1450
timestamp 1666464484
transform 1 0 163744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1454
timestamp 1666464484
transform 1 0 164192 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1457
timestamp 1666464484
transform 1 0 164528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1521
timestamp 1666464484
transform 1 0 171696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1525
timestamp 1666464484
transform 1 0 172144 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1528
timestamp 1666464484
transform 1 0 172480 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_1560
timestamp 1666464484
transform 1 0 176064 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1576
timestamp 1666464484
transform 1 0 177856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1580
timestamp 1666464484
transform 1 0 178304 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1666464484
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1666464484
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1666464484
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1666464484
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1666464484
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1666464484
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1666464484
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1666464484
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1666464484
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_215
timestamp 1666464484
transform 1 0 25424 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_247
timestamp 1666464484
transform 1 0 29008 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_263
timestamp 1666464484
transform 1 0 30800 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_277
timestamp 1666464484
transform 1 0 32368 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1666464484
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_286
timestamp 1666464484
transform 1 0 33376 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_302
timestamp 1666464484
transform 1 0 35168 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_306
timestamp 1666464484
transform 1 0 35616 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_310
timestamp 1666464484
transform 1 0 36064 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_314
timestamp 1666464484
transform 1 0 36512 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_316
timestamp 1666464484
transform 1 0 36736 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_319
timestamp 1666464484
transform 1 0 37072 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_323
timestamp 1666464484
transform 1 0 37520 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1666464484
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_357
timestamp 1666464484
transform 1 0 41328 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_360
timestamp 1666464484
transform 1 0 41664 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_364
timestamp 1666464484
transform 1 0 42112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_370
timestamp 1666464484
transform 1 0 42784 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_374
timestamp 1666464484
transform 1 0 43232 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_378
timestamp 1666464484
transform 1 0 43680 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_382
timestamp 1666464484
transform 1 0 44128 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_399
timestamp 1666464484
transform 1 0 46032 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_401
timestamp 1666464484
transform 1 0 46256 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_408
timestamp 1666464484
transform 1 0 47040 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1666464484
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1666464484
transform 1 0 49280 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_479
timestamp 1666464484
transform 1 0 54992 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_487
timestamp 1666464484
transform 1 0 55888 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_491
timestamp 1666464484
transform 1 0 56336 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_493
timestamp 1666464484
transform 1 0 56560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1666464484
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_499
timestamp 1666464484
transform 1 0 57232 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_518
timestamp 1666464484
transform 1 0 59360 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_522
timestamp 1666464484
transform 1 0 59808 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_526
timestamp 1666464484
transform 1 0 60256 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_556
timestamp 1666464484
transform 1 0 63616 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_558
timestamp 1666464484
transform 1 0 63840 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_565
timestamp 1666464484
transform 1 0 64624 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1666464484
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_570
timestamp 1666464484
transform 1 0 65184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_573
timestamp 1666464484
transform 1 0 65520 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_577
timestamp 1666464484
transform 1 0 65968 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_581
timestamp 1666464484
transform 1 0 66416 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_589
timestamp 1666464484
transform 1 0 67312 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_597
timestamp 1666464484
transform 1 0 68208 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_605
timestamp 1666464484
transform 1 0 69104 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1666464484
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_641
timestamp 1666464484
transform 1 0 73136 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_643
timestamp 1666464484
transform 1 0 73360 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_650
timestamp 1666464484
transform 1 0 74144 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_657
timestamp 1666464484
transform 1 0 74928 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_688
timestamp 1666464484
transform 1 0 78400 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_694
timestamp 1666464484
transform 1 0 79072 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_698
timestamp 1666464484
transform 1 0 79520 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_701
timestamp 1666464484
transform 1 0 79856 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_705
timestamp 1666464484
transform 1 0 80304 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1666464484
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_712
timestamp 1666464484
transform 1 0 81088 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_718
timestamp 1666464484
transform 1 0 81760 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_726
timestamp 1666464484
transform 1 0 82656 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_728
timestamp 1666464484
transform 1 0 82880 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_731
timestamp 1666464484
transform 1 0 83216 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_762
timestamp 1666464484
transform 1 0 86688 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_766
timestamp 1666464484
transform 1 0 87136 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_768
timestamp 1666464484
transform 1 0 87360 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_771
timestamp 1666464484
transform 1 0 87696 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_775
timestamp 1666464484
transform 1 0 88144 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_777
timestamp 1666464484
transform 1 0 88368 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1666464484
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_783
timestamp 1666464484
transform 1 0 89040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_789
timestamp 1666464484
transform 1 0 89712 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_822
timestamp 1666464484
transform 1 0 93408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_826
timestamp 1666464484
transform 1 0 93856 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_830
timestamp 1666464484
transform 1 0 94304 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_834
timestamp 1666464484
transform 1 0 94752 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_840
timestamp 1666464484
transform 1 0 95424 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1666464484
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_854
timestamp 1666464484
transform 1 0 96992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_859
timestamp 1666464484
transform 1 0 97552 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_873
timestamp 1666464484
transform 1 0 99120 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_883
timestamp 1666464484
transform 1 0 100240 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_887
timestamp 1666464484
transform 1 0 100688 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_891
timestamp 1666464484
transform 1 0 101136 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1666464484
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_925
timestamp 1666464484
transform 1 0 104944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_955
timestamp 1666464484
transform 1 0 108304 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_959
timestamp 1666464484
transform 1 0 108752 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_990
timestamp 1666464484
transform 1 0 112224 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_996
timestamp 1666464484
transform 1 0 112896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_999
timestamp 1666464484
transform 1 0 113232 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1003
timestamp 1666464484
transform 1 0 113680 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1007
timestamp 1666464484
transform 1 0 114128 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1011
timestamp 1666464484
transform 1 0 114576 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1015
timestamp 1666464484
transform 1 0 115024 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1023
timestamp 1666464484
transform 1 0 115920 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1031
timestamp 1666464484
transform 1 0 116816 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1039
timestamp 1666464484
transform 1 0 117712 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1043
timestamp 1666464484
transform 1 0 118160 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1050
timestamp 1666464484
transform 1 0 118944 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1054
timestamp 1666464484
transform 1 0 119392 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1058
timestamp 1666464484
transform 1 0 119840 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1062
timestamp 1666464484
transform 1 0 120288 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1064
timestamp 1666464484
transform 1 0 120512 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1067
timestamp 1666464484
transform 1 0 120848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1070
timestamp 1666464484
transform 1 0 121184 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1074
timestamp 1666464484
transform 1 0 121632 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_1078
timestamp 1666464484
transform 1 0 122080 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1110
timestamp 1666464484
transform 1 0 125664 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_1126
timestamp 1666464484
transform 1 0 127456 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1134
timestamp 1666464484
transform 1 0 128352 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1138
timestamp 1666464484
transform 1 0 128800 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1202
timestamp 1666464484
transform 1 0 135968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1206
timestamp 1666464484
transform 1 0 136416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1209
timestamp 1666464484
transform 1 0 136752 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1273
timestamp 1666464484
transform 1 0 143920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1277
timestamp 1666464484
transform 1 0 144368 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1280
timestamp 1666464484
transform 1 0 144704 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1344
timestamp 1666464484
transform 1 0 151872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1348
timestamp 1666464484
transform 1 0 152320 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1351
timestamp 1666464484
transform 1 0 152656 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1415
timestamp 1666464484
transform 1 0 159824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1419
timestamp 1666464484
transform 1 0 160272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1422
timestamp 1666464484
transform 1 0 160608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1486
timestamp 1666464484
transform 1 0 167776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1490
timestamp 1666464484
transform 1 0 168224 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1493
timestamp 1666464484
transform 1 0 168560 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1557
timestamp 1666464484
transform 1 0 175728 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1561
timestamp 1666464484
transform 1 0 176176 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1564
timestamp 1666464484
transform 1 0 176512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1580
timestamp 1666464484
transform 1 0 178304 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1666464484
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1666464484
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1666464484
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1666464484
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1666464484
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1666464484
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1666464484
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1666464484
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1666464484
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1666464484
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1666464484
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_250
timestamp 1666464484
transform 1 0 29344 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_258
timestamp 1666464484
transform 1 0 30240 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_289
timestamp 1666464484
transform 1 0 33712 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_293
timestamp 1666464484
transform 1 0 34160 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_301
timestamp 1666464484
transform 1 0 35056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_304
timestamp 1666464484
transform 1 0 35392 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_308
timestamp 1666464484
transform 1 0 35840 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_312
timestamp 1666464484
transform 1 0 36288 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_316
timestamp 1666464484
transform 1 0 36736 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1666464484
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_321
timestamp 1666464484
transform 1 0 37296 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_351
timestamp 1666464484
transform 1 0 40656 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_355
timestamp 1666464484
transform 1 0 41104 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_359
timestamp 1666464484
transform 1 0 41552 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_365
timestamp 1666464484
transform 1 0 42224 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_369
timestamp 1666464484
transform 1 0 42672 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_375
timestamp 1666464484
transform 1 0 43344 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_383
timestamp 1666464484
transform 1 0 44240 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1666464484
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1666464484
transform 1 0 45248 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_399
timestamp 1666464484
transform 1 0 46032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_432
timestamp 1666464484
transform 1 0 49728 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_440
timestamp 1666464484
transform 1 0 50624 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_444
timestamp 1666464484
transform 1 0 51072 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_452
timestamp 1666464484
transform 1 0 51968 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1666464484
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_463
timestamp 1666464484
transform 1 0 53200 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_469
timestamp 1666464484
transform 1 0 53872 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_486
timestamp 1666464484
transform 1 0 55776 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_517
timestamp 1666464484
transform 1 0 59248 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_519
timestamp 1666464484
transform 1 0 59472 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_522
timestamp 1666464484
transform 1 0 59808 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_530
timestamp 1666464484
transform 1 0 60704 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_534
timestamp 1666464484
transform 1 0 61152 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_540
timestamp 1666464484
transform 1 0 61824 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_544
timestamp 1666464484
transform 1 0 62272 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_548
timestamp 1666464484
transform 1 0 62720 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_552
timestamp 1666464484
transform 1 0 63168 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_556
timestamp 1666464484
transform 1 0 63616 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_560
timestamp 1666464484
transform 1 0 64064 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_564
timestamp 1666464484
transform 1 0 64512 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_568
timestamp 1666464484
transform 1 0 64960 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_601
timestamp 1666464484
transform 1 0 68656 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_605
timestamp 1666464484
transform 1 0 69104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_656
timestamp 1666464484
transform 1 0 74816 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_664
timestamp 1666464484
transform 1 0 75712 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_666
timestamp 1666464484
transform 1 0 75936 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1666464484
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_676
timestamp 1666464484
transform 1 0 77056 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_678
timestamp 1666464484
transform 1 0 77280 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_685
timestamp 1666464484
transform 1 0 78064 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_693
timestamp 1666464484
transform 1 0 78960 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_697
timestamp 1666464484
transform 1 0 79408 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_701
timestamp 1666464484
transform 1 0 79856 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_705
timestamp 1666464484
transform 1 0 80304 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_709
timestamp 1666464484
transform 1 0 80752 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_713
timestamp 1666464484
transform 1 0 81200 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_717
timestamp 1666464484
transform 1 0 81648 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_727
timestamp 1666464484
transform 1 0 82768 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_731
timestamp 1666464484
transform 1 0 83216 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_739
timestamp 1666464484
transform 1 0 84112 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_741
timestamp 1666464484
transform 1 0 84336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1666464484
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_747
timestamp 1666464484
transform 1 0 85008 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_749
timestamp 1666464484
transform 1 0 85232 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_752
timestamp 1666464484
transform 1 0 85568 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_756
timestamp 1666464484
transform 1 0 86016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_758
timestamp 1666464484
transform 1 0 86240 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_761
timestamp 1666464484
transform 1 0 86576 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_765
timestamp 1666464484
transform 1 0 87024 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_773
timestamp 1666464484
transform 1 0 87920 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_806
timestamp 1666464484
transform 1 0 91616 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_814
timestamp 1666464484
transform 1 0 92512 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_818
timestamp 1666464484
transform 1 0 92960 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_834
timestamp 1666464484
transform 1 0 94752 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_837
timestamp 1666464484
transform 1 0 95088 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_845
timestamp 1666464484
transform 1 0 95984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_855
timestamp 1666464484
transform 1 0 97104 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_868
timestamp 1666464484
transform 1 0 98560 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_877
timestamp 1666464484
transform 1 0 99568 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_881
timestamp 1666464484
transform 1 0 100016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_885
timestamp 1666464484
transform 1 0 100464 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_889
timestamp 1666464484
transform 1 0 100912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_892
timestamp 1666464484
transform 1 0 101248 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_896
timestamp 1666464484
transform 1 0 101696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_900
timestamp 1666464484
transform 1 0 102144 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_907
timestamp 1666464484
transform 1 0 102928 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_911
timestamp 1666464484
transform 1 0 103376 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_915
timestamp 1666464484
transform 1 0 103824 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_919
timestamp 1666464484
transform 1 0 104272 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_921
timestamp 1666464484
transform 1 0 104496 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_924
timestamp 1666464484
transform 1 0 104832 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_928
timestamp 1666464484
transform 1 0 105280 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_932
timestamp 1666464484
transform 1 0 105728 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_936
timestamp 1666464484
transform 1 0 106176 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_940
timestamp 1666464484
transform 1 0 106624 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_944
timestamp 1666464484
transform 1 0 107072 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_948
timestamp 1666464484
transform 1 0 107520 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_950
timestamp 1666464484
transform 1 0 107744 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_953
timestamp 1666464484
transform 1 0 108080 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1666464484
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_960
timestamp 1666464484
transform 1 0 108864 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_993
timestamp 1666464484
transform 1 0 112560 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_997
timestamp 1666464484
transform 1 0 113008 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1001
timestamp 1666464484
transform 1 0 113456 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1005
timestamp 1666464484
transform 1 0 113904 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1009
timestamp 1666464484
transform 1 0 114352 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1013
timestamp 1666464484
transform 1 0 114800 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1017
timestamp 1666464484
transform 1 0 115248 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1021
timestamp 1666464484
transform 1 0 115696 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1025
timestamp 1666464484
transform 1 0 116144 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1031
timestamp 1666464484
transform 1 0 116816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1038
timestamp 1666464484
transform 1 0 117600 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1048
timestamp 1666464484
transform 1 0 118720 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1056
timestamp 1666464484
transform 1 0 119616 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_1060
timestamp 1666464484
transform 1 0 120064 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_1092
timestamp 1666464484
transform 1 0 123648 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1102
timestamp 1666464484
transform 1 0 124768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1166
timestamp 1666464484
transform 1 0 131936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1170
timestamp 1666464484
transform 1 0 132384 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1173
timestamp 1666464484
transform 1 0 132720 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1237
timestamp 1666464484
transform 1 0 139888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1241
timestamp 1666464484
transform 1 0 140336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1244
timestamp 1666464484
transform 1 0 140672 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1308
timestamp 1666464484
transform 1 0 147840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1312
timestamp 1666464484
transform 1 0 148288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1315
timestamp 1666464484
transform 1 0 148624 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1379
timestamp 1666464484
transform 1 0 155792 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1383
timestamp 1666464484
transform 1 0 156240 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1386
timestamp 1666464484
transform 1 0 156576 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1450
timestamp 1666464484
transform 1 0 163744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1454
timestamp 1666464484
transform 1 0 164192 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1457
timestamp 1666464484
transform 1 0 164528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1521
timestamp 1666464484
transform 1 0 171696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1525
timestamp 1666464484
transform 1 0 172144 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_1528
timestamp 1666464484
transform 1 0 172480 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_1560
timestamp 1666464484
transform 1 0 176064 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1576
timestamp 1666464484
transform 1 0 177856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1580
timestamp 1666464484
transform 1 0 178304 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1666464484
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1666464484
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1666464484
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1666464484
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1666464484
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1666464484
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1666464484
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1666464484
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1666464484
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1666464484
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1666464484
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_286
timestamp 1666464484
transform 1 0 33376 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_318
timestamp 1666464484
transform 1 0 36960 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_322
timestamp 1666464484
transform 1 0 37408 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_329
timestamp 1666464484
transform 1 0 38192 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_333
timestamp 1666464484
transform 1 0 38640 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_336
timestamp 1666464484
transform 1 0 38976 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_338
timestamp 1666464484
transform 1 0 39200 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_341
timestamp 1666464484
transform 1 0 39536 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_345
timestamp 1666464484
transform 1 0 39984 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_353
timestamp 1666464484
transform 1 0 40880 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_357
timestamp 1666464484
transform 1 0 41328 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_365
timestamp 1666464484
transform 1 0 42224 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_396
timestamp 1666464484
transform 1 0 45696 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_400
timestamp 1666464484
transform 1 0 46144 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_404
timestamp 1666464484
transform 1 0 46592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_410
timestamp 1666464484
transform 1 0 47264 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_418
timestamp 1666464484
transform 1 0 48160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_422
timestamp 1666464484
transform 1 0 48608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1666464484
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_428
timestamp 1666464484
transform 1 0 49280 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_434
timestamp 1666464484
transform 1 0 49952 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_438
timestamp 1666464484
transform 1 0 50400 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_442
timestamp 1666464484
transform 1 0 50848 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_446
timestamp 1666464484
transform 1 0 51296 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_452
timestamp 1666464484
transform 1 0 51968 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_454
timestamp 1666464484
transform 1 0 52192 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_484
timestamp 1666464484
transform 1 0 55552 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_490
timestamp 1666464484
transform 1 0 56224 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_494
timestamp 1666464484
transform 1 0 56672 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1666464484
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_499
timestamp 1666464484
transform 1 0 57232 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_506
timestamp 1666464484
transform 1 0 58016 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_510
timestamp 1666464484
transform 1 0 58464 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_514
timestamp 1666464484
transform 1 0 58912 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_547
timestamp 1666464484
transform 1 0 62608 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_551
timestamp 1666464484
transform 1 0 63056 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_555
timestamp 1666464484
transform 1 0 63504 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_559
timestamp 1666464484
transform 1 0 63952 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_563
timestamp 1666464484
transform 1 0 64400 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1666464484
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_570
timestamp 1666464484
transform 1 0 65184 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_574
timestamp 1666464484
transform 1 0 65632 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_605
timestamp 1666464484
transform 1 0 69104 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1666464484
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_641
timestamp 1666464484
transform 1 0 73136 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_645
timestamp 1666464484
transform 1 0 73584 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_653
timestamp 1666464484
transform 1 0 74480 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_660
timestamp 1666464484
transform 1 0 75264 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_666
timestamp 1666464484
transform 1 0 75936 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_670
timestamp 1666464484
transform 1 0 76384 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_703
timestamp 1666464484
transform 1 0 80080 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_705
timestamp 1666464484
transform 1 0 80304 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_708
timestamp 1666464484
transform 1 0 80640 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_712
timestamp 1666464484
transform 1 0 81088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_715
timestamp 1666464484
transform 1 0 81424 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_723
timestamp 1666464484
transform 1 0 82320 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_754
timestamp 1666464484
transform 1 0 85792 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_762
timestamp 1666464484
transform 1 0 86688 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_766
timestamp 1666464484
transform 1 0 87136 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_772
timestamp 1666464484
transform 1 0 87808 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1666464484
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_783
timestamp 1666464484
transform 1 0 89040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_815
timestamp 1666464484
transform 1 0 92624 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_831
timestamp 1666464484
transform 1 0 94416 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_839
timestamp 1666464484
transform 1 0 95312 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_843
timestamp 1666464484
transform 1 0 95760 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_847
timestamp 1666464484
transform 1 0 96208 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1666464484
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_854
timestamp 1666464484
transform 1 0 96992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_884
timestamp 1666464484
transform 1 0 100352 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_888
timestamp 1666464484
transform 1 0 100800 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_892
timestamp 1666464484
transform 1 0 101248 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_896
timestamp 1666464484
transform 1 0 101696 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_900
timestamp 1666464484
transform 1 0 102144 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_904
timestamp 1666464484
transform 1 0 102592 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_908
timestamp 1666464484
transform 1 0 103040 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_914
timestamp 1666464484
transform 1 0 103712 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1666464484
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_925
timestamp 1666464484
transform 1 0 104944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_932
timestamp 1666464484
transform 1 0 105728 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_936
timestamp 1666464484
transform 1 0 106176 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_940
timestamp 1666464484
transform 1 0 106624 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_944
timestamp 1666464484
transform 1 0 107072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_948
timestamp 1666464484
transform 1 0 107520 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_952
timestamp 1666464484
transform 1 0 107968 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_955
timestamp 1666464484
transform 1 0 108304 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_959
timestamp 1666464484
transform 1 0 108752 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_992
timestamp 1666464484
transform 1 0 112448 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_996
timestamp 1666464484
transform 1 0 112896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_999
timestamp 1666464484
transform 1 0 113232 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1003
timestamp 1666464484
transform 1 0 113680 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1007
timestamp 1666464484
transform 1 0 114128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1011
timestamp 1666464484
transform 1 0 114576 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1013
timestamp 1666464484
transform 1 0 114800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1016
timestamp 1666464484
transform 1 0 115136 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1020
timestamp 1666464484
transform 1 0 115584 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1024
timestamp 1666464484
transform 1 0 116032 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1028
timestamp 1666464484
transform 1 0 116480 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1032
timestamp 1666464484
transform 1 0 116928 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1036
timestamp 1666464484
transform 1 0 117376 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1040
timestamp 1666464484
transform 1 0 117824 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_1044
timestamp 1666464484
transform 1 0 118272 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1060
timestamp 1666464484
transform 1 0 120064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1064
timestamp 1666464484
transform 1 0 120512 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1067
timestamp 1666464484
transform 1 0 120848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1131
timestamp 1666464484
transform 1 0 128016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1135
timestamp 1666464484
transform 1 0 128464 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1138
timestamp 1666464484
transform 1 0 128800 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1202
timestamp 1666464484
transform 1 0 135968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1206
timestamp 1666464484
transform 1 0 136416 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1209
timestamp 1666464484
transform 1 0 136752 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1273
timestamp 1666464484
transform 1 0 143920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1277
timestamp 1666464484
transform 1 0 144368 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1280
timestamp 1666464484
transform 1 0 144704 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1344
timestamp 1666464484
transform 1 0 151872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1348
timestamp 1666464484
transform 1 0 152320 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1351
timestamp 1666464484
transform 1 0 152656 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1415
timestamp 1666464484
transform 1 0 159824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1419
timestamp 1666464484
transform 1 0 160272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1422
timestamp 1666464484
transform 1 0 160608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1486
timestamp 1666464484
transform 1 0 167776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1490
timestamp 1666464484
transform 1 0 168224 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1493
timestamp 1666464484
transform 1 0 168560 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1557
timestamp 1666464484
transform 1 0 175728 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1561
timestamp 1666464484
transform 1 0 176176 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_1564
timestamp 1666464484
transform 1 0 176512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1580
timestamp 1666464484
transform 1 0 178304 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1666464484
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1666464484
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1666464484
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1666464484
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1666464484
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1666464484
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1666464484
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1666464484
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1666464484
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1666464484
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1666464484
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1666464484
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1666464484
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1666464484
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_321
timestamp 1666464484
transform 1 0 37296 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_329
timestamp 1666464484
transform 1 0 38192 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_333
timestamp 1666464484
transform 1 0 38640 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_335
timestamp 1666464484
transform 1 0 38864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_338
timestamp 1666464484
transform 1 0 39200 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_342
timestamp 1666464484
transform 1 0 39648 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_374
timestamp 1666464484
transform 1 0 43232 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_392
timestamp 1666464484
transform 1 0 45248 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_400
timestamp 1666464484
transform 1 0 46144 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_402
timestamp 1666464484
transform 1 0 46368 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_405
timestamp 1666464484
transform 1 0 46704 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_407
timestamp 1666464484
transform 1 0 46928 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_410
timestamp 1666464484
transform 1 0 47264 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_414
timestamp 1666464484
transform 1 0 47712 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_418
timestamp 1666464484
transform 1 0 48160 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_424
timestamp 1666464484
transform 1 0 48832 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_440
timestamp 1666464484
transform 1 0 50624 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_446
timestamp 1666464484
transform 1 0 51296 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_450
timestamp 1666464484
transform 1 0 51744 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_454
timestamp 1666464484
transform 1 0 52192 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1666464484
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_463
timestamp 1666464484
transform 1 0 53200 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_465
timestamp 1666464484
transform 1 0 53424 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_472
timestamp 1666464484
transform 1 0 54208 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_476
timestamp 1666464484
transform 1 0 54656 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_478
timestamp 1666464484
transform 1 0 54880 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_481
timestamp 1666464484
transform 1 0 55216 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_485
timestamp 1666464484
transform 1 0 55664 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_489
timestamp 1666464484
transform 1 0 56112 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_493
timestamp 1666464484
transform 1 0 56560 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_497
timestamp 1666464484
transform 1 0 57008 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_499
timestamp 1666464484
transform 1 0 57232 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_502
timestamp 1666464484
transform 1 0 57568 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_506
timestamp 1666464484
transform 1 0 58016 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_510
timestamp 1666464484
transform 1 0 58464 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_514
timestamp 1666464484
transform 1 0 58912 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_524
timestamp 1666464484
transform 1 0 60032 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_528
timestamp 1666464484
transform 1 0 60480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_534
timestamp 1666464484
transform 1 0 61152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_537
timestamp 1666464484
transform 1 0 61488 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_541
timestamp 1666464484
transform 1 0 61936 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_545
timestamp 1666464484
transform 1 0 62384 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_549
timestamp 1666464484
transform 1 0 62832 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_553
timestamp 1666464484
transform 1 0 63280 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_555
timestamp 1666464484
transform 1 0 63504 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_585
timestamp 1666464484
transform 1 0 66864 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_589
timestamp 1666464484
transform 1 0 67312 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_591
timestamp 1666464484
transform 1 0 67536 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_594
timestamp 1666464484
transform 1 0 67872 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_598
timestamp 1666464484
transform 1 0 68320 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1666464484
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_605
timestamp 1666464484
transform 1 0 69104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_608
timestamp 1666464484
transform 1 0 69440 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_612
timestamp 1666464484
transform 1 0 69888 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_616
timestamp 1666464484
transform 1 0 70336 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_623
timestamp 1666464484
transform 1 0 71120 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_631
timestamp 1666464484
transform 1 0 72016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_666
timestamp 1666464484
transform 1 0 75936 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_670
timestamp 1666464484
transform 1 0 76384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_676
timestamp 1666464484
transform 1 0 77056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_679
timestamp 1666464484
transform 1 0 77392 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_683
timestamp 1666464484
transform 1 0 77840 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_686
timestamp 1666464484
transform 1 0 78176 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_690
timestamp 1666464484
transform 1 0 78624 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_694
timestamp 1666464484
transform 1 0 79072 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_725
timestamp 1666464484
transform 1 0 82544 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_729
timestamp 1666464484
transform 1 0 82992 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_737
timestamp 1666464484
transform 1 0 83888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_741
timestamp 1666464484
transform 1 0 84336 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1666464484
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_747
timestamp 1666464484
transform 1 0 85008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_779
timestamp 1666464484
transform 1 0 88592 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_781
timestamp 1666464484
transform 1 0 88816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_784
timestamp 1666464484
transform 1 0 89152 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1666464484
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_818
timestamp 1666464484
transform 1 0 92960 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_822
timestamp 1666464484
transform 1 0 93408 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_824
timestamp 1666464484
transform 1 0 93632 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_827
timestamp 1666464484
transform 1 0 93968 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_858
timestamp 1666464484
transform 1 0 97440 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_862
timestamp 1666464484
transform 1 0 97888 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_866
timestamp 1666464484
transform 1 0 98336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_870
timestamp 1666464484
transform 1 0 98784 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_877
timestamp 1666464484
transform 1 0 99568 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_881
timestamp 1666464484
transform 1 0 100016 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_885
timestamp 1666464484
transform 1 0 100464 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_889
timestamp 1666464484
transform 1 0 100912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_892
timestamp 1666464484
transform 1 0 101248 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_896
timestamp 1666464484
transform 1 0 101696 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_900
timestamp 1666464484
transform 1 0 102144 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_904
timestamp 1666464484
transform 1 0 102592 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_908
timestamp 1666464484
transform 1 0 103040 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_941
timestamp 1666464484
transform 1 0 106736 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_945
timestamp 1666464484
transform 1 0 107184 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_949
timestamp 1666464484
transform 1 0 107632 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_953
timestamp 1666464484
transform 1 0 108080 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_957
timestamp 1666464484
transform 1 0 108528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_960
timestamp 1666464484
transform 1 0 108864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_992
timestamp 1666464484
transform 1 0 112448 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_996
timestamp 1666464484
transform 1 0 112896 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_1000
timestamp 1666464484
transform 1 0 113344 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1008
timestamp 1666464484
transform 1 0 114240 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1010
timestamp 1666464484
transform 1 0 114464 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1013
timestamp 1666464484
transform 1 0 114800 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1015
timestamp 1666464484
transform 1 0 115024 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_1018
timestamp 1666464484
transform 1 0 115360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1026
timestamp 1666464484
transform 1 0 116256 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1666464484
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1031
timestamp 1666464484
transform 1 0 116816 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1095
timestamp 1666464484
transform 1 0 123984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1099
timestamp 1666464484
transform 1 0 124432 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1102
timestamp 1666464484
transform 1 0 124768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1166
timestamp 1666464484
transform 1 0 131936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1170
timestamp 1666464484
transform 1 0 132384 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1173
timestamp 1666464484
transform 1 0 132720 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1237
timestamp 1666464484
transform 1 0 139888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1241
timestamp 1666464484
transform 1 0 140336 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1244
timestamp 1666464484
transform 1 0 140672 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1308
timestamp 1666464484
transform 1 0 147840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1312
timestamp 1666464484
transform 1 0 148288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1315
timestamp 1666464484
transform 1 0 148624 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1379
timestamp 1666464484
transform 1 0 155792 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1383
timestamp 1666464484
transform 1 0 156240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1386
timestamp 1666464484
transform 1 0 156576 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1450
timestamp 1666464484
transform 1 0 163744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1454
timestamp 1666464484
transform 1 0 164192 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1457
timestamp 1666464484
transform 1 0 164528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1521
timestamp 1666464484
transform 1 0 171696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1525
timestamp 1666464484
transform 1 0 172144 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_1528
timestamp 1666464484
transform 1 0 172480 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_1560
timestamp 1666464484
transform 1 0 176064 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1576
timestamp 1666464484
transform 1 0 177856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1580
timestamp 1666464484
transform 1 0 178304 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1666464484
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1666464484
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1666464484
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1666464484
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1666464484
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1666464484
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1666464484
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1666464484
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1666464484
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1666464484
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1666464484
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1666464484
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1666464484
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1666464484
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1666464484
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1666464484
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1666464484
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1666464484
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_428
timestamp 1666464484
transform 1 0 49280 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_444
timestamp 1666464484
transform 1 0 51072 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_452
timestamp 1666464484
transform 1 0 51968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_456
timestamp 1666464484
transform 1 0 52416 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_460
timestamp 1666464484
transform 1 0 52864 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_476
timestamp 1666464484
transform 1 0 54656 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_478
timestamp 1666464484
transform 1 0 54880 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_481
timestamp 1666464484
transform 1 0 55216 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_499
timestamp 1666464484
transform 1 0 57232 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_502
timestamp 1666464484
transform 1 0 57568 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_506
timestamp 1666464484
transform 1 0 58016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_510
timestamp 1666464484
transform 1 0 58464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_514
timestamp 1666464484
transform 1 0 58912 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_518
timestamp 1666464484
transform 1 0 59360 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_522
timestamp 1666464484
transform 1 0 59808 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_539
timestamp 1666464484
transform 1 0 61712 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_543
timestamp 1666464484
transform 1 0 62160 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_551
timestamp 1666464484
transform 1 0 63056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_555
timestamp 1666464484
transform 1 0 63504 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_559
timestamp 1666464484
transform 1 0 63952 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_563
timestamp 1666464484
transform 1 0 64400 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1666464484
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_570
timestamp 1666464484
transform 1 0 65184 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_576
timestamp 1666464484
transform 1 0 65856 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_580
timestamp 1666464484
transform 1 0 66304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_584
timestamp 1666464484
transform 1 0 66752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_587
timestamp 1666464484
transform 1 0 67088 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_591
timestamp 1666464484
transform 1 0 67536 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_595
timestamp 1666464484
transform 1 0 67984 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_598
timestamp 1666464484
transform 1 0 68320 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_602
timestamp 1666464484
transform 1 0 68768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_606
timestamp 1666464484
transform 1 0 69216 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_610
timestamp 1666464484
transform 1 0 69664 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_616
timestamp 1666464484
transform 1 0 70336 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_620
timestamp 1666464484
transform 1 0 70784 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_624
timestamp 1666464484
transform 1 0 71232 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_628
timestamp 1666464484
transform 1 0 71680 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_631
timestamp 1666464484
transform 1 0 72016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_635
timestamp 1666464484
transform 1 0 72464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_641
timestamp 1666464484
transform 1 0 73136 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_647
timestamp 1666464484
transform 1 0 73808 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_651
timestamp 1666464484
transform 1 0 74256 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_655
timestamp 1666464484
transform 1 0 74704 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_659
timestamp 1666464484
transform 1 0 75152 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_663
timestamp 1666464484
transform 1 0 75600 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_669
timestamp 1666464484
transform 1 0 76272 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_673
timestamp 1666464484
transform 1 0 76720 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_677
timestamp 1666464484
transform 1 0 77168 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_681
timestamp 1666464484
transform 1 0 77616 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_685
timestamp 1666464484
transform 1 0 78064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_691
timestamp 1666464484
transform 1 0 78736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_697
timestamp 1666464484
transform 1 0 79408 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_701
timestamp 1666464484
transform 1 0 79856 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_705
timestamp 1666464484
transform 1 0 80304 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1666464484
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_712
timestamp 1666464484
transform 1 0 81088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_715
timestamp 1666464484
transform 1 0 81424 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_719
timestamp 1666464484
transform 1 0 81872 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_723
timestamp 1666464484
transform 1 0 82320 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_727
timestamp 1666464484
transform 1 0 82768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_729
timestamp 1666464484
transform 1 0 82992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_732
timestamp 1666464484
transform 1 0 83328 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_736
timestamp 1666464484
transform 1 0 83776 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_740
timestamp 1666464484
transform 1 0 84224 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_746
timestamp 1666464484
transform 1 0 84896 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_756
timestamp 1666464484
transform 1 0 86016 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_772
timestamp 1666464484
transform 1 0 87808 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1666464484
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_783
timestamp 1666464484
transform 1 0 89040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_791
timestamp 1666464484
transform 1 0 89936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_797
timestamp 1666464484
transform 1 0 90608 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_805
timestamp 1666464484
transform 1 0 91504 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_837
timestamp 1666464484
transform 1 0 95088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_845
timestamp 1666464484
transform 1 0 95984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_849
timestamp 1666464484
transform 1 0 96432 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1666464484
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_854
timestamp 1666464484
transform 1 0 96992 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_862
timestamp 1666464484
transform 1 0 97888 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_866
timestamp 1666464484
transform 1 0 98336 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_899
timestamp 1666464484
transform 1 0 102032 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_915
timestamp 1666464484
transform 1 0 103824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_919
timestamp 1666464484
transform 1 0 104272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_922
timestamp 1666464484
transform 1 0 104608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_925
timestamp 1666464484
transform 1 0 104944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_955
timestamp 1666464484
transform 1 0 108304 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_986
timestamp 1666464484
transform 1 0 111776 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_990
timestamp 1666464484
transform 1 0 112224 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_996
timestamp 1666464484
transform 1 0 112896 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1060
timestamp 1666464484
transform 1 0 120064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1064
timestamp 1666464484
transform 1 0 120512 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1067
timestamp 1666464484
transform 1 0 120848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1131
timestamp 1666464484
transform 1 0 128016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1135
timestamp 1666464484
transform 1 0 128464 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1138
timestamp 1666464484
transform 1 0 128800 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1202
timestamp 1666464484
transform 1 0 135968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1206
timestamp 1666464484
transform 1 0 136416 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1209
timestamp 1666464484
transform 1 0 136752 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1273
timestamp 1666464484
transform 1 0 143920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1277
timestamp 1666464484
transform 1 0 144368 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1280
timestamp 1666464484
transform 1 0 144704 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1344
timestamp 1666464484
transform 1 0 151872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1348
timestamp 1666464484
transform 1 0 152320 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1351
timestamp 1666464484
transform 1 0 152656 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1415
timestamp 1666464484
transform 1 0 159824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1419
timestamp 1666464484
transform 1 0 160272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1422
timestamp 1666464484
transform 1 0 160608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1486
timestamp 1666464484
transform 1 0 167776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1490
timestamp 1666464484
transform 1 0 168224 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1493
timestamp 1666464484
transform 1 0 168560 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1557
timestamp 1666464484
transform 1 0 175728 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1561
timestamp 1666464484
transform 1 0 176176 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_1564
timestamp 1666464484
transform 1 0 176512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1580
timestamp 1666464484
transform 1 0 178304 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1666464484
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1666464484
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1666464484
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1666464484
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1666464484
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1666464484
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1666464484
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1666464484
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1666464484
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1666464484
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1666464484
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1666464484
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1666464484
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1666464484
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1666464484
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1666464484
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1666464484
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1666464484
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1666464484
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1666464484
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1666464484
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1666464484
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_534
timestamp 1666464484
transform 1 0 61152 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_566
timestamp 1666464484
transform 1 0 64736 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_582
timestamp 1666464484
transform 1 0 66528 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_586
timestamp 1666464484
transform 1 0 66976 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_588
timestamp 1666464484
transform 1 0 67200 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_591
timestamp 1666464484
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_595
timestamp 1666464484
transform 1 0 67984 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_598
timestamp 1666464484
transform 1 0 68320 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1666464484
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_605
timestamp 1666464484
transform 1 0 69104 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_611
timestamp 1666464484
transform 1 0 69776 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_615
timestamp 1666464484
transform 1 0 70224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_621
timestamp 1666464484
transform 1 0 70896 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_625
timestamp 1666464484
transform 1 0 71344 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_629
timestamp 1666464484
transform 1 0 71792 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_631
timestamp 1666464484
transform 1 0 72016 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_634
timestamp 1666464484
transform 1 0 72352 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_638
timestamp 1666464484
transform 1 0 72800 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_642
timestamp 1666464484
transform 1 0 73248 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_646
timestamp 1666464484
transform 1 0 73696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_652
timestamp 1666464484
transform 1 0 74368 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_656
timestamp 1666464484
transform 1 0 74816 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_660
timestamp 1666464484
transform 1 0 75264 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_662
timestamp 1666464484
transform 1 0 75488 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_665
timestamp 1666464484
transform 1 0 75824 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_669
timestamp 1666464484
transform 1 0 76272 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1666464484
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_676
timestamp 1666464484
transform 1 0 77056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_679
timestamp 1666464484
transform 1 0 77392 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_683
timestamp 1666464484
transform 1 0 77840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_687
timestamp 1666464484
transform 1 0 78288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_690
timestamp 1666464484
transform 1 0 78624 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_692
timestamp 1666464484
transform 1 0 78848 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_695
timestamp 1666464484
transform 1 0 79184 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_697
timestamp 1666464484
transform 1 0 79408 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_700
timestamp 1666464484
transform 1 0 79744 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_704
timestamp 1666464484
transform 1 0 80192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_708
timestamp 1666464484
transform 1 0 80640 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_711
timestamp 1666464484
transform 1 0 80976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_717
timestamp 1666464484
transform 1 0 81648 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_727
timestamp 1666464484
transform 1 0 82768 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_731
timestamp 1666464484
transform 1 0 83216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_739
timestamp 1666464484
transform 1 0 84112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_743
timestamp 1666464484
transform 1 0 84560 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1666464484
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1666464484
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1666464484
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1666464484
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_882
timestamp 1666464484
transform 1 0 100128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1666464484
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_889
timestamp 1666464484
transform 1 0 100912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_919
timestamp 1666464484
transform 1 0 104272 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_951
timestamp 1666464484
transform 1 0 107856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_955
timestamp 1666464484
transform 1 0 108304 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_957
timestamp 1666464484
transform 1 0 108528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1666464484
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1666464484
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1666464484
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1031
timestamp 1666464484
transform 1 0 116816 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1095
timestamp 1666464484
transform 1 0 123984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1099
timestamp 1666464484
transform 1 0 124432 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1102
timestamp 1666464484
transform 1 0 124768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1166
timestamp 1666464484
transform 1 0 131936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1170
timestamp 1666464484
transform 1 0 132384 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1173
timestamp 1666464484
transform 1 0 132720 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1237
timestamp 1666464484
transform 1 0 139888 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1241
timestamp 1666464484
transform 1 0 140336 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1244
timestamp 1666464484
transform 1 0 140672 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1308
timestamp 1666464484
transform 1 0 147840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1312
timestamp 1666464484
transform 1 0 148288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1315
timestamp 1666464484
transform 1 0 148624 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1379
timestamp 1666464484
transform 1 0 155792 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1383
timestamp 1666464484
transform 1 0 156240 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1386
timestamp 1666464484
transform 1 0 156576 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1450
timestamp 1666464484
transform 1 0 163744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1454
timestamp 1666464484
transform 1 0 164192 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1457
timestamp 1666464484
transform 1 0 164528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1521
timestamp 1666464484
transform 1 0 171696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1525
timestamp 1666464484
transform 1 0 172144 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_1528
timestamp 1666464484
transform 1 0 172480 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_1560
timestamp 1666464484
transform 1 0 176064 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1576
timestamp 1666464484
transform 1 0 177856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1580
timestamp 1666464484
transform 1 0 178304 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1666464484
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1666464484
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1666464484
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1666464484
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1666464484
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1666464484
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1666464484
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1666464484
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1666464484
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1666464484
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1666464484
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1666464484
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1666464484
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1666464484
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1666464484
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1666464484
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1666464484
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1666464484
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1666464484
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1666464484
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1666464484
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1666464484
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1666464484
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1666464484
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_570
timestamp 1666464484
transform 1 0 65184 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_602
timestamp 1666464484
transform 1 0 68768 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_606
timestamp 1666464484
transform 1 0 69216 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_610
timestamp 1666464484
transform 1 0 69664 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_612
timestamp 1666464484
transform 1 0 69888 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_615
timestamp 1666464484
transform 1 0 70224 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_619
timestamp 1666464484
transform 1 0 70672 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_623
timestamp 1666464484
transform 1 0 71120 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_631
timestamp 1666464484
transform 1 0 72016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_635
timestamp 1666464484
transform 1 0 72464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1666464484
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_641
timestamp 1666464484
transform 1 0 73136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_649
timestamp 1666464484
transform 1 0 74032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_653
timestamp 1666464484
transform 1 0 74480 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_655
timestamp 1666464484
transform 1 0 74704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_658
timestamp 1666464484
transform 1 0 75040 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_660
timestamp 1666464484
transform 1 0 75264 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_663
timestamp 1666464484
transform 1 0 75600 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_667
timestamp 1666464484
transform 1 0 76048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_677
timestamp 1666464484
transform 1 0 77168 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_687
timestamp 1666464484
transform 1 0 78288 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_691
timestamp 1666464484
transform 1 0 78736 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_695
timestamp 1666464484
transform 1 0 79184 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_701
timestamp 1666464484
transform 1 0 79856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_705
timestamp 1666464484
transform 1 0 80304 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1666464484
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1666464484
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1666464484
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1666464484
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1666464484
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1666464484
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1666464484
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1666464484
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1666464484
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1666464484
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1666464484
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1666464484
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1666464484
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_996
timestamp 1666464484
transform 1 0 112896 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1060
timestamp 1666464484
transform 1 0 120064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1064
timestamp 1666464484
transform 1 0 120512 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1067
timestamp 1666464484
transform 1 0 120848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1131
timestamp 1666464484
transform 1 0 128016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1135
timestamp 1666464484
transform 1 0 128464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1138
timestamp 1666464484
transform 1 0 128800 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1202
timestamp 1666464484
transform 1 0 135968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1206
timestamp 1666464484
transform 1 0 136416 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1209
timestamp 1666464484
transform 1 0 136752 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1273
timestamp 1666464484
transform 1 0 143920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1277
timestamp 1666464484
transform 1 0 144368 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1280
timestamp 1666464484
transform 1 0 144704 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1344
timestamp 1666464484
transform 1 0 151872 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1348
timestamp 1666464484
transform 1 0 152320 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1351
timestamp 1666464484
transform 1 0 152656 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1415
timestamp 1666464484
transform 1 0 159824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1419
timestamp 1666464484
transform 1 0 160272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1422
timestamp 1666464484
transform 1 0 160608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1486
timestamp 1666464484
transform 1 0 167776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1490
timestamp 1666464484
transform 1 0 168224 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1493
timestamp 1666464484
transform 1 0 168560 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1557
timestamp 1666464484
transform 1 0 175728 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1561
timestamp 1666464484
transform 1 0 176176 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_1564
timestamp 1666464484
transform 1 0 176512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1580
timestamp 1666464484
transform 1 0 178304 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1666464484
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1666464484
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1666464484
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1666464484
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1666464484
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1666464484
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1666464484
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1666464484
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1666464484
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1666464484
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1666464484
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1666464484
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1666464484
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1666464484
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1666464484
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1666464484
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1666464484
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1666464484
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1666464484
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1666464484
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1666464484
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1666464484
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1666464484
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1666464484
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1666464484
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1666464484
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1666464484
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1666464484
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1666464484
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1666464484
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1666464484
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1666464484
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1666464484
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1666464484
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1666464484
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1666464484
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1666464484
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1666464484
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1666464484
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1666464484
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_960
timestamp 1666464484
transform 1 0 108864 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1024
timestamp 1666464484
transform 1 0 116032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1028
timestamp 1666464484
transform 1 0 116480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1031
timestamp 1666464484
transform 1 0 116816 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1095
timestamp 1666464484
transform 1 0 123984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1099
timestamp 1666464484
transform 1 0 124432 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1102
timestamp 1666464484
transform 1 0 124768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1166
timestamp 1666464484
transform 1 0 131936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1170
timestamp 1666464484
transform 1 0 132384 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1173
timestamp 1666464484
transform 1 0 132720 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1237
timestamp 1666464484
transform 1 0 139888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1241
timestamp 1666464484
transform 1 0 140336 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1244
timestamp 1666464484
transform 1 0 140672 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1308
timestamp 1666464484
transform 1 0 147840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1312
timestamp 1666464484
transform 1 0 148288 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1315
timestamp 1666464484
transform 1 0 148624 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1379
timestamp 1666464484
transform 1 0 155792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1383
timestamp 1666464484
transform 1 0 156240 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1386
timestamp 1666464484
transform 1 0 156576 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1450
timestamp 1666464484
transform 1 0 163744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1454
timestamp 1666464484
transform 1 0 164192 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1457
timestamp 1666464484
transform 1 0 164528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1521
timestamp 1666464484
transform 1 0 171696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1525
timestamp 1666464484
transform 1 0 172144 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_1528
timestamp 1666464484
transform 1 0 172480 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_1560
timestamp 1666464484
transform 1 0 176064 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1576
timestamp 1666464484
transform 1 0 177856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1580
timestamp 1666464484
transform 1 0 178304 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1666464484
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1666464484
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1666464484
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1666464484
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1666464484
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1666464484
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1666464484
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1666464484
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1666464484
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1666464484
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1666464484
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1666464484
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1666464484
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1666464484
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1666464484
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1666464484
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1666464484
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1666464484
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1666464484
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1666464484
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1666464484
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1666464484
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1666464484
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1666464484
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1666464484
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1666464484
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1666464484
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1666464484
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1666464484
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1666464484
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1666464484
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1666464484
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1666464484
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1666464484
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1666464484
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1666464484
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1666464484
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1666464484
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1666464484
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1666464484
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1666464484
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1666464484
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_996
timestamp 1666464484
transform 1 0 112896 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1060
timestamp 1666464484
transform 1 0 120064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1064
timestamp 1666464484
transform 1 0 120512 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1067
timestamp 1666464484
transform 1 0 120848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1131
timestamp 1666464484
transform 1 0 128016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1135
timestamp 1666464484
transform 1 0 128464 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1138
timestamp 1666464484
transform 1 0 128800 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1202
timestamp 1666464484
transform 1 0 135968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1206
timestamp 1666464484
transform 1 0 136416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1209
timestamp 1666464484
transform 1 0 136752 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1273
timestamp 1666464484
transform 1 0 143920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1277
timestamp 1666464484
transform 1 0 144368 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1280
timestamp 1666464484
transform 1 0 144704 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1344
timestamp 1666464484
transform 1 0 151872 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1348
timestamp 1666464484
transform 1 0 152320 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1351
timestamp 1666464484
transform 1 0 152656 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1415
timestamp 1666464484
transform 1 0 159824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1419
timestamp 1666464484
transform 1 0 160272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1422
timestamp 1666464484
transform 1 0 160608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1486
timestamp 1666464484
transform 1 0 167776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1490
timestamp 1666464484
transform 1 0 168224 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1493
timestamp 1666464484
transform 1 0 168560 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1557
timestamp 1666464484
transform 1 0 175728 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1561
timestamp 1666464484
transform 1 0 176176 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_1564
timestamp 1666464484
transform 1 0 176512 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1580
timestamp 1666464484
transform 1 0 178304 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1666464484
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1666464484
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1666464484
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1666464484
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1666464484
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1666464484
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1666464484
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1666464484
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1666464484
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1666464484
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1666464484
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1666464484
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1666464484
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1666464484
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1666464484
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1666464484
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1666464484
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1666464484
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1666464484
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1666464484
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1666464484
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1666464484
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1666464484
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1666464484
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1666464484
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1666464484
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1666464484
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1666464484
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_676
timestamp 1666464484
transform 1 0 77056 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_740
timestamp 1666464484
transform 1 0 84224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_744
timestamp 1666464484
transform 1 0 84672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_747
timestamp 1666464484
transform 1 0 85008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_811
timestamp 1666464484
transform 1 0 92176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_815
timestamp 1666464484
transform 1 0 92624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_818
timestamp 1666464484
transform 1 0 92960 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_882
timestamp 1666464484
transform 1 0 100128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_886
timestamp 1666464484
transform 1 0 100576 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_889
timestamp 1666464484
transform 1 0 100912 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_953
timestamp 1666464484
transform 1 0 108080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_957
timestamp 1666464484
transform 1 0 108528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_960
timestamp 1666464484
transform 1 0 108864 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1024
timestamp 1666464484
transform 1 0 116032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1028
timestamp 1666464484
transform 1 0 116480 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1031
timestamp 1666464484
transform 1 0 116816 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1095
timestamp 1666464484
transform 1 0 123984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1099
timestamp 1666464484
transform 1 0 124432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1102
timestamp 1666464484
transform 1 0 124768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1166
timestamp 1666464484
transform 1 0 131936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1170
timestamp 1666464484
transform 1 0 132384 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1173
timestamp 1666464484
transform 1 0 132720 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1237
timestamp 1666464484
transform 1 0 139888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1241
timestamp 1666464484
transform 1 0 140336 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1244
timestamp 1666464484
transform 1 0 140672 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1308
timestamp 1666464484
transform 1 0 147840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1312
timestamp 1666464484
transform 1 0 148288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1315
timestamp 1666464484
transform 1 0 148624 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1379
timestamp 1666464484
transform 1 0 155792 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1383
timestamp 1666464484
transform 1 0 156240 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1386
timestamp 1666464484
transform 1 0 156576 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1450
timestamp 1666464484
transform 1 0 163744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1454
timestamp 1666464484
transform 1 0 164192 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1457
timestamp 1666464484
transform 1 0 164528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1521
timestamp 1666464484
transform 1 0 171696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1525
timestamp 1666464484
transform 1 0 172144 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_1528
timestamp 1666464484
transform 1 0 172480 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1560
timestamp 1666464484
transform 1 0 176064 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1576
timestamp 1666464484
transform 1 0 177856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1580
timestamp 1666464484
transform 1 0 178304 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1666464484
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1666464484
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1666464484
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1666464484
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1666464484
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1666464484
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1666464484
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1666464484
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1666464484
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1666464484
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1666464484
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1666464484
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1666464484
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1666464484
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1666464484
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1666464484
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1666464484
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1666464484
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1666464484
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1666464484
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1666464484
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1666464484
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1666464484
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1666464484
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1666464484
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1666464484
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1666464484
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_641
timestamp 1666464484
transform 1 0 73136 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_705
timestamp 1666464484
transform 1 0 80304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_709
timestamp 1666464484
transform 1 0 80752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_712
timestamp 1666464484
transform 1 0 81088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_776
timestamp 1666464484
transform 1 0 88256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_780
timestamp 1666464484
transform 1 0 88704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_783
timestamp 1666464484
transform 1 0 89040 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_847
timestamp 1666464484
transform 1 0 96208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_851
timestamp 1666464484
transform 1 0 96656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_854
timestamp 1666464484
transform 1 0 96992 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_918
timestamp 1666464484
transform 1 0 104160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_922
timestamp 1666464484
transform 1 0 104608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_925
timestamp 1666464484
transform 1 0 104944 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_989
timestamp 1666464484
transform 1 0 112112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_993
timestamp 1666464484
transform 1 0 112560 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_996
timestamp 1666464484
transform 1 0 112896 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1060
timestamp 1666464484
transform 1 0 120064 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1064
timestamp 1666464484
transform 1 0 120512 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1067
timestamp 1666464484
transform 1 0 120848 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1131
timestamp 1666464484
transform 1 0 128016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1135
timestamp 1666464484
transform 1 0 128464 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1138
timestamp 1666464484
transform 1 0 128800 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1202
timestamp 1666464484
transform 1 0 135968 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1206
timestamp 1666464484
transform 1 0 136416 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1209
timestamp 1666464484
transform 1 0 136752 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1273
timestamp 1666464484
transform 1 0 143920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1277
timestamp 1666464484
transform 1 0 144368 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1280
timestamp 1666464484
transform 1 0 144704 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1344
timestamp 1666464484
transform 1 0 151872 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1348
timestamp 1666464484
transform 1 0 152320 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1351
timestamp 1666464484
transform 1 0 152656 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1415
timestamp 1666464484
transform 1 0 159824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1419
timestamp 1666464484
transform 1 0 160272 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1422
timestamp 1666464484
transform 1 0 160608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1486
timestamp 1666464484
transform 1 0 167776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1490
timestamp 1666464484
transform 1 0 168224 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1493
timestamp 1666464484
transform 1 0 168560 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1557
timestamp 1666464484
transform 1 0 175728 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1561
timestamp 1666464484
transform 1 0 176176 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_1564
timestamp 1666464484
transform 1 0 176512 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1580
timestamp 1666464484
transform 1 0 178304 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1666464484
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1666464484
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1666464484
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1666464484
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1666464484
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1666464484
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1666464484
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1666464484
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1666464484
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1666464484
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1666464484
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1666464484
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1666464484
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1666464484
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1666464484
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1666464484
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1666464484
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1666464484
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1666464484
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1666464484
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1666464484
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1666464484
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1666464484
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1666464484
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1666464484
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1666464484
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1666464484
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1666464484
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_676
timestamp 1666464484
transform 1 0 77056 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_740
timestamp 1666464484
transform 1 0 84224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_744
timestamp 1666464484
transform 1 0 84672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_747
timestamp 1666464484
transform 1 0 85008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_811
timestamp 1666464484
transform 1 0 92176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_815
timestamp 1666464484
transform 1 0 92624 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_818
timestamp 1666464484
transform 1 0 92960 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_882
timestamp 1666464484
transform 1 0 100128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_886
timestamp 1666464484
transform 1 0 100576 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_889
timestamp 1666464484
transform 1 0 100912 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_953
timestamp 1666464484
transform 1 0 108080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_957
timestamp 1666464484
transform 1 0 108528 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_960
timestamp 1666464484
transform 1 0 108864 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1024
timestamp 1666464484
transform 1 0 116032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1028
timestamp 1666464484
transform 1 0 116480 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1031
timestamp 1666464484
transform 1 0 116816 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1095
timestamp 1666464484
transform 1 0 123984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1099
timestamp 1666464484
transform 1 0 124432 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1102
timestamp 1666464484
transform 1 0 124768 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1166
timestamp 1666464484
transform 1 0 131936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1170
timestamp 1666464484
transform 1 0 132384 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1173
timestamp 1666464484
transform 1 0 132720 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1237
timestamp 1666464484
transform 1 0 139888 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1241
timestamp 1666464484
transform 1 0 140336 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1244
timestamp 1666464484
transform 1 0 140672 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1308
timestamp 1666464484
transform 1 0 147840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1312
timestamp 1666464484
transform 1 0 148288 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1315
timestamp 1666464484
transform 1 0 148624 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1379
timestamp 1666464484
transform 1 0 155792 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1383
timestamp 1666464484
transform 1 0 156240 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1386
timestamp 1666464484
transform 1 0 156576 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1450
timestamp 1666464484
transform 1 0 163744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1454
timestamp 1666464484
transform 1 0 164192 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1457
timestamp 1666464484
transform 1 0 164528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1521
timestamp 1666464484
transform 1 0 171696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1525
timestamp 1666464484
transform 1 0 172144 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_1528
timestamp 1666464484
transform 1 0 172480 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_1560
timestamp 1666464484
transform 1 0 176064 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1576
timestamp 1666464484
transform 1 0 177856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1580
timestamp 1666464484
transform 1 0 178304 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1666464484
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1666464484
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1666464484
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1666464484
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1666464484
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1666464484
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1666464484
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1666464484
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1666464484
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1666464484
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1666464484
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1666464484
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1666464484
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1666464484
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1666464484
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1666464484
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1666464484
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1666464484
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1666464484
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1666464484
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1666464484
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1666464484
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1666464484
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1666464484
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1666464484
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1666464484
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1666464484
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_641
timestamp 1666464484
transform 1 0 73136 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_705
timestamp 1666464484
transform 1 0 80304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_709
timestamp 1666464484
transform 1 0 80752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_712
timestamp 1666464484
transform 1 0 81088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_776
timestamp 1666464484
transform 1 0 88256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_780
timestamp 1666464484
transform 1 0 88704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_783
timestamp 1666464484
transform 1 0 89040 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_847
timestamp 1666464484
transform 1 0 96208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_851
timestamp 1666464484
transform 1 0 96656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_854
timestamp 1666464484
transform 1 0 96992 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_918
timestamp 1666464484
transform 1 0 104160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_922
timestamp 1666464484
transform 1 0 104608 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_925
timestamp 1666464484
transform 1 0 104944 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_989
timestamp 1666464484
transform 1 0 112112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_993
timestamp 1666464484
transform 1 0 112560 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_996
timestamp 1666464484
transform 1 0 112896 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1060
timestamp 1666464484
transform 1 0 120064 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1064
timestamp 1666464484
transform 1 0 120512 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1067
timestamp 1666464484
transform 1 0 120848 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1131
timestamp 1666464484
transform 1 0 128016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1135
timestamp 1666464484
transform 1 0 128464 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1138
timestamp 1666464484
transform 1 0 128800 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1202
timestamp 1666464484
transform 1 0 135968 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1206
timestamp 1666464484
transform 1 0 136416 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1209
timestamp 1666464484
transform 1 0 136752 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1273
timestamp 1666464484
transform 1 0 143920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1277
timestamp 1666464484
transform 1 0 144368 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1280
timestamp 1666464484
transform 1 0 144704 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1344
timestamp 1666464484
transform 1 0 151872 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1348
timestamp 1666464484
transform 1 0 152320 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1351
timestamp 1666464484
transform 1 0 152656 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1415
timestamp 1666464484
transform 1 0 159824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1419
timestamp 1666464484
transform 1 0 160272 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1422
timestamp 1666464484
transform 1 0 160608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1486
timestamp 1666464484
transform 1 0 167776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1490
timestamp 1666464484
transform 1 0 168224 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1493
timestamp 1666464484
transform 1 0 168560 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1557
timestamp 1666464484
transform 1 0 175728 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1561
timestamp 1666464484
transform 1 0 176176 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_1564
timestamp 1666464484
transform 1 0 176512 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1580
timestamp 1666464484
transform 1 0 178304 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1666464484
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1666464484
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1666464484
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1666464484
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1666464484
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1666464484
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1666464484
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1666464484
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1666464484
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1666464484
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1666464484
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1666464484
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1666464484
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1666464484
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1666464484
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1666464484
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1666464484
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1666464484
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1666464484
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1666464484
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1666464484
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1666464484
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1666464484
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1666464484
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1666464484
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1666464484
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1666464484
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_676
timestamp 1666464484
transform 1 0 77056 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_740
timestamp 1666464484
transform 1 0 84224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_744
timestamp 1666464484
transform 1 0 84672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_747
timestamp 1666464484
transform 1 0 85008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_811
timestamp 1666464484
transform 1 0 92176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_815
timestamp 1666464484
transform 1 0 92624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_818
timestamp 1666464484
transform 1 0 92960 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_882
timestamp 1666464484
transform 1 0 100128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_886
timestamp 1666464484
transform 1 0 100576 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_889
timestamp 1666464484
transform 1 0 100912 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_953
timestamp 1666464484
transform 1 0 108080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_957
timestamp 1666464484
transform 1 0 108528 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_960
timestamp 1666464484
transform 1 0 108864 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1024
timestamp 1666464484
transform 1 0 116032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1028
timestamp 1666464484
transform 1 0 116480 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1031
timestamp 1666464484
transform 1 0 116816 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1095
timestamp 1666464484
transform 1 0 123984 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1099
timestamp 1666464484
transform 1 0 124432 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1102
timestamp 1666464484
transform 1 0 124768 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1166
timestamp 1666464484
transform 1 0 131936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1170
timestamp 1666464484
transform 1 0 132384 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1173
timestamp 1666464484
transform 1 0 132720 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1237
timestamp 1666464484
transform 1 0 139888 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1241
timestamp 1666464484
transform 1 0 140336 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1244
timestamp 1666464484
transform 1 0 140672 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1308
timestamp 1666464484
transform 1 0 147840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1312
timestamp 1666464484
transform 1 0 148288 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1315
timestamp 1666464484
transform 1 0 148624 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1379
timestamp 1666464484
transform 1 0 155792 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1383
timestamp 1666464484
transform 1 0 156240 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1386
timestamp 1666464484
transform 1 0 156576 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1450
timestamp 1666464484
transform 1 0 163744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1454
timestamp 1666464484
transform 1 0 164192 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1457
timestamp 1666464484
transform 1 0 164528 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1521
timestamp 1666464484
transform 1 0 171696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1525
timestamp 1666464484
transform 1 0 172144 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_1528
timestamp 1666464484
transform 1 0 172480 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_1560
timestamp 1666464484
transform 1 0 176064 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1576
timestamp 1666464484
transform 1 0 177856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1580
timestamp 1666464484
transform 1 0 178304 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1666464484
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1666464484
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1666464484
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1666464484
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1666464484
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1666464484
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1666464484
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1666464484
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1666464484
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1666464484
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1666464484
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1666464484
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1666464484
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1666464484
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1666464484
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1666464484
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1666464484
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1666464484
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1666464484
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1666464484
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1666464484
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1666464484
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1666464484
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1666464484
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1666464484
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1666464484
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_641
timestamp 1666464484
transform 1 0 73136 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_705
timestamp 1666464484
transform 1 0 80304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_709
timestamp 1666464484
transform 1 0 80752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_712
timestamp 1666464484
transform 1 0 81088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_776
timestamp 1666464484
transform 1 0 88256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_780
timestamp 1666464484
transform 1 0 88704 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_783
timestamp 1666464484
transform 1 0 89040 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_847
timestamp 1666464484
transform 1 0 96208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_851
timestamp 1666464484
transform 1 0 96656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_854
timestamp 1666464484
transform 1 0 96992 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_918
timestamp 1666464484
transform 1 0 104160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_922
timestamp 1666464484
transform 1 0 104608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_925
timestamp 1666464484
transform 1 0 104944 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_989
timestamp 1666464484
transform 1 0 112112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_993
timestamp 1666464484
transform 1 0 112560 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_996
timestamp 1666464484
transform 1 0 112896 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1060
timestamp 1666464484
transform 1 0 120064 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1064
timestamp 1666464484
transform 1 0 120512 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1067
timestamp 1666464484
transform 1 0 120848 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1131
timestamp 1666464484
transform 1 0 128016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1135
timestamp 1666464484
transform 1 0 128464 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1138
timestamp 1666464484
transform 1 0 128800 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1202
timestamp 1666464484
transform 1 0 135968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1206
timestamp 1666464484
transform 1 0 136416 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1209
timestamp 1666464484
transform 1 0 136752 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1273
timestamp 1666464484
transform 1 0 143920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1277
timestamp 1666464484
transform 1 0 144368 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1280
timestamp 1666464484
transform 1 0 144704 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1344
timestamp 1666464484
transform 1 0 151872 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1348
timestamp 1666464484
transform 1 0 152320 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1351
timestamp 1666464484
transform 1 0 152656 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1415
timestamp 1666464484
transform 1 0 159824 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1419
timestamp 1666464484
transform 1 0 160272 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1422
timestamp 1666464484
transform 1 0 160608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1486
timestamp 1666464484
transform 1 0 167776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1490
timestamp 1666464484
transform 1 0 168224 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1493
timestamp 1666464484
transform 1 0 168560 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1557
timestamp 1666464484
transform 1 0 175728 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1561
timestamp 1666464484
transform 1 0 176176 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_1564
timestamp 1666464484
transform 1 0 176512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1580
timestamp 1666464484
transform 1 0 178304 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1666464484
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1666464484
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1666464484
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1666464484
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1666464484
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1666464484
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1666464484
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1666464484
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1666464484
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1666464484
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1666464484
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1666464484
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1666464484
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1666464484
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1666464484
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1666464484
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1666464484
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1666464484
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1666464484
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1666464484
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1666464484
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1666464484
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1666464484
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1666464484
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1666464484
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1666464484
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1666464484
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1666464484
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_676
timestamp 1666464484
transform 1 0 77056 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_740
timestamp 1666464484
transform 1 0 84224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_744
timestamp 1666464484
transform 1 0 84672 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_747
timestamp 1666464484
transform 1 0 85008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_811
timestamp 1666464484
transform 1 0 92176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_815
timestamp 1666464484
transform 1 0 92624 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_818
timestamp 1666464484
transform 1 0 92960 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_882
timestamp 1666464484
transform 1 0 100128 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_886
timestamp 1666464484
transform 1 0 100576 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_889
timestamp 1666464484
transform 1 0 100912 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_953
timestamp 1666464484
transform 1 0 108080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_957
timestamp 1666464484
transform 1 0 108528 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_960
timestamp 1666464484
transform 1 0 108864 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1024
timestamp 1666464484
transform 1 0 116032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1028
timestamp 1666464484
transform 1 0 116480 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1031
timestamp 1666464484
transform 1 0 116816 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1095
timestamp 1666464484
transform 1 0 123984 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1099
timestamp 1666464484
transform 1 0 124432 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1102
timestamp 1666464484
transform 1 0 124768 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1166
timestamp 1666464484
transform 1 0 131936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1170
timestamp 1666464484
transform 1 0 132384 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1173
timestamp 1666464484
transform 1 0 132720 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1237
timestamp 1666464484
transform 1 0 139888 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1241
timestamp 1666464484
transform 1 0 140336 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1244
timestamp 1666464484
transform 1 0 140672 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1308
timestamp 1666464484
transform 1 0 147840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1312
timestamp 1666464484
transform 1 0 148288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1315
timestamp 1666464484
transform 1 0 148624 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1379
timestamp 1666464484
transform 1 0 155792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1383
timestamp 1666464484
transform 1 0 156240 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1386
timestamp 1666464484
transform 1 0 156576 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1450
timestamp 1666464484
transform 1 0 163744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1454
timestamp 1666464484
transform 1 0 164192 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1457
timestamp 1666464484
transform 1 0 164528 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1521
timestamp 1666464484
transform 1 0 171696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1525
timestamp 1666464484
transform 1 0 172144 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_1528
timestamp 1666464484
transform 1 0 172480 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_1560
timestamp 1666464484
transform 1 0 176064 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1576
timestamp 1666464484
transform 1 0 177856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1580
timestamp 1666464484
transform 1 0 178304 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1666464484
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1666464484
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1666464484
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1666464484
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1666464484
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1666464484
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1666464484
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1666464484
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1666464484
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1666464484
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1666464484
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1666464484
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1666464484
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1666464484
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1666464484
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1666464484
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1666464484
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1666464484
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1666464484
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1666464484
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1666464484
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1666464484
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1666464484
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1666464484
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1666464484
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1666464484
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1666464484
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_641
timestamp 1666464484
transform 1 0 73136 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_705
timestamp 1666464484
transform 1 0 80304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_709
timestamp 1666464484
transform 1 0 80752 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_712
timestamp 1666464484
transform 1 0 81088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_776
timestamp 1666464484
transform 1 0 88256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_780
timestamp 1666464484
transform 1 0 88704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_783
timestamp 1666464484
transform 1 0 89040 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_847
timestamp 1666464484
transform 1 0 96208 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_851
timestamp 1666464484
transform 1 0 96656 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_854
timestamp 1666464484
transform 1 0 96992 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_918
timestamp 1666464484
transform 1 0 104160 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_922
timestamp 1666464484
transform 1 0 104608 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_925
timestamp 1666464484
transform 1 0 104944 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_989
timestamp 1666464484
transform 1 0 112112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_993
timestamp 1666464484
transform 1 0 112560 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_996
timestamp 1666464484
transform 1 0 112896 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1060
timestamp 1666464484
transform 1 0 120064 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1064
timestamp 1666464484
transform 1 0 120512 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1067
timestamp 1666464484
transform 1 0 120848 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1131
timestamp 1666464484
transform 1 0 128016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1135
timestamp 1666464484
transform 1 0 128464 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1138
timestamp 1666464484
transform 1 0 128800 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1202
timestamp 1666464484
transform 1 0 135968 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1206
timestamp 1666464484
transform 1 0 136416 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1209
timestamp 1666464484
transform 1 0 136752 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1273
timestamp 1666464484
transform 1 0 143920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1277
timestamp 1666464484
transform 1 0 144368 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1280
timestamp 1666464484
transform 1 0 144704 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1344
timestamp 1666464484
transform 1 0 151872 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1348
timestamp 1666464484
transform 1 0 152320 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1351
timestamp 1666464484
transform 1 0 152656 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1415
timestamp 1666464484
transform 1 0 159824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1419
timestamp 1666464484
transform 1 0 160272 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1422
timestamp 1666464484
transform 1 0 160608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1486
timestamp 1666464484
transform 1 0 167776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1490
timestamp 1666464484
transform 1 0 168224 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1493
timestamp 1666464484
transform 1 0 168560 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1557
timestamp 1666464484
transform 1 0 175728 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1561
timestamp 1666464484
transform 1 0 176176 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_1564
timestamp 1666464484
transform 1 0 176512 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1580
timestamp 1666464484
transform 1 0 178304 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1666464484
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1666464484
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1666464484
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1666464484
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1666464484
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1666464484
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1666464484
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1666464484
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1666464484
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1666464484
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1666464484
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1666464484
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1666464484
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1666464484
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1666464484
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1666464484
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1666464484
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1666464484
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1666464484
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1666464484
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1666464484
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1666464484
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1666464484
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1666464484
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1666464484
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1666464484
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1666464484
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_669
timestamp 1666464484
transform 1 0 76272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1666464484
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_676
timestamp 1666464484
transform 1 0 77056 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_740
timestamp 1666464484
transform 1 0 84224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_744
timestamp 1666464484
transform 1 0 84672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_747
timestamp 1666464484
transform 1 0 85008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_811
timestamp 1666464484
transform 1 0 92176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_815
timestamp 1666464484
transform 1 0 92624 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_818
timestamp 1666464484
transform 1 0 92960 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_882
timestamp 1666464484
transform 1 0 100128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_886
timestamp 1666464484
transform 1 0 100576 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_889
timestamp 1666464484
transform 1 0 100912 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_953
timestamp 1666464484
transform 1 0 108080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_957
timestamp 1666464484
transform 1 0 108528 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_960
timestamp 1666464484
transform 1 0 108864 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1024
timestamp 1666464484
transform 1 0 116032 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1028
timestamp 1666464484
transform 1 0 116480 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1031
timestamp 1666464484
transform 1 0 116816 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1095
timestamp 1666464484
transform 1 0 123984 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1099
timestamp 1666464484
transform 1 0 124432 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1102
timestamp 1666464484
transform 1 0 124768 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1166
timestamp 1666464484
transform 1 0 131936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1170
timestamp 1666464484
transform 1 0 132384 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1173
timestamp 1666464484
transform 1 0 132720 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1237
timestamp 1666464484
transform 1 0 139888 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1241
timestamp 1666464484
transform 1 0 140336 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1244
timestamp 1666464484
transform 1 0 140672 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1308
timestamp 1666464484
transform 1 0 147840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1312
timestamp 1666464484
transform 1 0 148288 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1315
timestamp 1666464484
transform 1 0 148624 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1379
timestamp 1666464484
transform 1 0 155792 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1383
timestamp 1666464484
transform 1 0 156240 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1386
timestamp 1666464484
transform 1 0 156576 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1450
timestamp 1666464484
transform 1 0 163744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1454
timestamp 1666464484
transform 1 0 164192 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1457
timestamp 1666464484
transform 1 0 164528 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1521
timestamp 1666464484
transform 1 0 171696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1525
timestamp 1666464484
transform 1 0 172144 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_1528
timestamp 1666464484
transform 1 0 172480 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_1560
timestamp 1666464484
transform 1 0 176064 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1576
timestamp 1666464484
transform 1 0 177856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1580
timestamp 1666464484
transform 1 0 178304 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1666464484
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1666464484
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1666464484
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1666464484
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1666464484
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1666464484
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1666464484
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1666464484
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1666464484
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1666464484
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1666464484
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1666464484
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1666464484
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1666464484
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1666464484
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1666464484
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1666464484
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1666464484
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1666464484
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1666464484
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1666464484
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1666464484
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1666464484
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1666464484
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1666464484
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1666464484
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1666464484
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_641
timestamp 1666464484
transform 1 0 73136 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_705
timestamp 1666464484
transform 1 0 80304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_709
timestamp 1666464484
transform 1 0 80752 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_712
timestamp 1666464484
transform 1 0 81088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_776
timestamp 1666464484
transform 1 0 88256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_780
timestamp 1666464484
transform 1 0 88704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_783
timestamp 1666464484
transform 1 0 89040 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_847
timestamp 1666464484
transform 1 0 96208 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_851
timestamp 1666464484
transform 1 0 96656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_854
timestamp 1666464484
transform 1 0 96992 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_918
timestamp 1666464484
transform 1 0 104160 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_922
timestamp 1666464484
transform 1 0 104608 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_925
timestamp 1666464484
transform 1 0 104944 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_989
timestamp 1666464484
transform 1 0 112112 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_993
timestamp 1666464484
transform 1 0 112560 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_996
timestamp 1666464484
transform 1 0 112896 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1060
timestamp 1666464484
transform 1 0 120064 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1064
timestamp 1666464484
transform 1 0 120512 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1067
timestamp 1666464484
transform 1 0 120848 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1131
timestamp 1666464484
transform 1 0 128016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1135
timestamp 1666464484
transform 1 0 128464 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1138
timestamp 1666464484
transform 1 0 128800 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1202
timestamp 1666464484
transform 1 0 135968 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1206
timestamp 1666464484
transform 1 0 136416 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1209
timestamp 1666464484
transform 1 0 136752 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1273
timestamp 1666464484
transform 1 0 143920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1277
timestamp 1666464484
transform 1 0 144368 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1280
timestamp 1666464484
transform 1 0 144704 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1344
timestamp 1666464484
transform 1 0 151872 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1348
timestamp 1666464484
transform 1 0 152320 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1351
timestamp 1666464484
transform 1 0 152656 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1415
timestamp 1666464484
transform 1 0 159824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1419
timestamp 1666464484
transform 1 0 160272 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1422
timestamp 1666464484
transform 1 0 160608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1486
timestamp 1666464484
transform 1 0 167776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1490
timestamp 1666464484
transform 1 0 168224 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1493
timestamp 1666464484
transform 1 0 168560 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1557
timestamp 1666464484
transform 1 0 175728 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1561
timestamp 1666464484
transform 1 0 176176 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_1564
timestamp 1666464484
transform 1 0 176512 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1580
timestamp 1666464484
transform 1 0 178304 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1666464484
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1666464484
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1666464484
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1666464484
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1666464484
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1666464484
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1666464484
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1666464484
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1666464484
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1666464484
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1666464484
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1666464484
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1666464484
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1666464484
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1666464484
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1666464484
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1666464484
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1666464484
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1666464484
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1666464484
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1666464484
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1666464484
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1666464484
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1666464484
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1666464484
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1666464484
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1666464484
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1666464484
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_676
timestamp 1666464484
transform 1 0 77056 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_740
timestamp 1666464484
transform 1 0 84224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_744
timestamp 1666464484
transform 1 0 84672 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_747
timestamp 1666464484
transform 1 0 85008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_811
timestamp 1666464484
transform 1 0 92176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_815
timestamp 1666464484
transform 1 0 92624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_818
timestamp 1666464484
transform 1 0 92960 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_882
timestamp 1666464484
transform 1 0 100128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_886
timestamp 1666464484
transform 1 0 100576 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_889
timestamp 1666464484
transform 1 0 100912 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_953
timestamp 1666464484
transform 1 0 108080 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_957
timestamp 1666464484
transform 1 0 108528 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_960
timestamp 1666464484
transform 1 0 108864 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1024
timestamp 1666464484
transform 1 0 116032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1028
timestamp 1666464484
transform 1 0 116480 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1031
timestamp 1666464484
transform 1 0 116816 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1095
timestamp 1666464484
transform 1 0 123984 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1099
timestamp 1666464484
transform 1 0 124432 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1102
timestamp 1666464484
transform 1 0 124768 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1166
timestamp 1666464484
transform 1 0 131936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1170
timestamp 1666464484
transform 1 0 132384 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1173
timestamp 1666464484
transform 1 0 132720 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1237
timestamp 1666464484
transform 1 0 139888 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1241
timestamp 1666464484
transform 1 0 140336 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1244
timestamp 1666464484
transform 1 0 140672 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1308
timestamp 1666464484
transform 1 0 147840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1312
timestamp 1666464484
transform 1 0 148288 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1315
timestamp 1666464484
transform 1 0 148624 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1379
timestamp 1666464484
transform 1 0 155792 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1383
timestamp 1666464484
transform 1 0 156240 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1386
timestamp 1666464484
transform 1 0 156576 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1450
timestamp 1666464484
transform 1 0 163744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1454
timestamp 1666464484
transform 1 0 164192 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1457
timestamp 1666464484
transform 1 0 164528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1521
timestamp 1666464484
transform 1 0 171696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1525
timestamp 1666464484
transform 1 0 172144 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_1528
timestamp 1666464484
transform 1 0 172480 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_1560
timestamp 1666464484
transform 1 0 176064 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1576
timestamp 1666464484
transform 1 0 177856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1580
timestamp 1666464484
transform 1 0 178304 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1666464484
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1666464484
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1666464484
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1666464484
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1666464484
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1666464484
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1666464484
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1666464484
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1666464484
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1666464484
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1666464484
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1666464484
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1666464484
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1666464484
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1666464484
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1666464484
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1666464484
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1666464484
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1666464484
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1666464484
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1666464484
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1666464484
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1666464484
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1666464484
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1666464484
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1666464484
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1666464484
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_641
timestamp 1666464484
transform 1 0 73136 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_705
timestamp 1666464484
transform 1 0 80304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_709
timestamp 1666464484
transform 1 0 80752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_712
timestamp 1666464484
transform 1 0 81088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_776
timestamp 1666464484
transform 1 0 88256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_780
timestamp 1666464484
transform 1 0 88704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_783
timestamp 1666464484
transform 1 0 89040 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_847
timestamp 1666464484
transform 1 0 96208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_851
timestamp 1666464484
transform 1 0 96656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_854
timestamp 1666464484
transform 1 0 96992 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_918
timestamp 1666464484
transform 1 0 104160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_922
timestamp 1666464484
transform 1 0 104608 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_925
timestamp 1666464484
transform 1 0 104944 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_989
timestamp 1666464484
transform 1 0 112112 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_993
timestamp 1666464484
transform 1 0 112560 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_996
timestamp 1666464484
transform 1 0 112896 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1060
timestamp 1666464484
transform 1 0 120064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1064
timestamp 1666464484
transform 1 0 120512 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1067
timestamp 1666464484
transform 1 0 120848 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1131
timestamp 1666464484
transform 1 0 128016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1135
timestamp 1666464484
transform 1 0 128464 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1138
timestamp 1666464484
transform 1 0 128800 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1202
timestamp 1666464484
transform 1 0 135968 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1206
timestamp 1666464484
transform 1 0 136416 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1209
timestamp 1666464484
transform 1 0 136752 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1273
timestamp 1666464484
transform 1 0 143920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1277
timestamp 1666464484
transform 1 0 144368 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1280
timestamp 1666464484
transform 1 0 144704 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1344
timestamp 1666464484
transform 1 0 151872 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1348
timestamp 1666464484
transform 1 0 152320 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1351
timestamp 1666464484
transform 1 0 152656 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1415
timestamp 1666464484
transform 1 0 159824 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1419
timestamp 1666464484
transform 1 0 160272 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1422
timestamp 1666464484
transform 1 0 160608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1486
timestamp 1666464484
transform 1 0 167776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1490
timestamp 1666464484
transform 1 0 168224 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1493
timestamp 1666464484
transform 1 0 168560 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1557
timestamp 1666464484
transform 1 0 175728 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1561
timestamp 1666464484
transform 1 0 176176 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_1564
timestamp 1666464484
transform 1 0 176512 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1580
timestamp 1666464484
transform 1 0 178304 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1666464484
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1666464484
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1666464484
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1666464484
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1666464484
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1666464484
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1666464484
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1666464484
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1666464484
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1666464484
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1666464484
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1666464484
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1666464484
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1666464484
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1666464484
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1666464484
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1666464484
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1666464484
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1666464484
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1666464484
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1666464484
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1666464484
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1666464484
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1666464484
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1666464484
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1666464484
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1666464484
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1666464484
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_676
timestamp 1666464484
transform 1 0 77056 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_740
timestamp 1666464484
transform 1 0 84224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_744
timestamp 1666464484
transform 1 0 84672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_747
timestamp 1666464484
transform 1 0 85008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_811
timestamp 1666464484
transform 1 0 92176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_815
timestamp 1666464484
transform 1 0 92624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_818
timestamp 1666464484
transform 1 0 92960 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_882
timestamp 1666464484
transform 1 0 100128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_886
timestamp 1666464484
transform 1 0 100576 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_889
timestamp 1666464484
transform 1 0 100912 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_953
timestamp 1666464484
transform 1 0 108080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_957
timestamp 1666464484
transform 1 0 108528 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_960
timestamp 1666464484
transform 1 0 108864 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1024
timestamp 1666464484
transform 1 0 116032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1028
timestamp 1666464484
transform 1 0 116480 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1031
timestamp 1666464484
transform 1 0 116816 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1095
timestamp 1666464484
transform 1 0 123984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1099
timestamp 1666464484
transform 1 0 124432 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1102
timestamp 1666464484
transform 1 0 124768 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1166
timestamp 1666464484
transform 1 0 131936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1170
timestamp 1666464484
transform 1 0 132384 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1173
timestamp 1666464484
transform 1 0 132720 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1237
timestamp 1666464484
transform 1 0 139888 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1241
timestamp 1666464484
transform 1 0 140336 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1244
timestamp 1666464484
transform 1 0 140672 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1308
timestamp 1666464484
transform 1 0 147840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1312
timestamp 1666464484
transform 1 0 148288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1315
timestamp 1666464484
transform 1 0 148624 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1379
timestamp 1666464484
transform 1 0 155792 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1383
timestamp 1666464484
transform 1 0 156240 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1386
timestamp 1666464484
transform 1 0 156576 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1450
timestamp 1666464484
transform 1 0 163744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1454
timestamp 1666464484
transform 1 0 164192 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1457
timestamp 1666464484
transform 1 0 164528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1521
timestamp 1666464484
transform 1 0 171696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1525
timestamp 1666464484
transform 1 0 172144 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_1528
timestamp 1666464484
transform 1 0 172480 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_1560
timestamp 1666464484
transform 1 0 176064 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1576
timestamp 1666464484
transform 1 0 177856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1580
timestamp 1666464484
transform 1 0 178304 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1666464484
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1666464484
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1666464484
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1666464484
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1666464484
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1666464484
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1666464484
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1666464484
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1666464484
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1666464484
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1666464484
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1666464484
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1666464484
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1666464484
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1666464484
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1666464484
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1666464484
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1666464484
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1666464484
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1666464484
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1666464484
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1666464484
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1666464484
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1666464484
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1666464484
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1666464484
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_641
timestamp 1666464484
transform 1 0 73136 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_705
timestamp 1666464484
transform 1 0 80304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_709
timestamp 1666464484
transform 1 0 80752 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_712
timestamp 1666464484
transform 1 0 81088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_776
timestamp 1666464484
transform 1 0 88256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_780
timestamp 1666464484
transform 1 0 88704 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_783
timestamp 1666464484
transform 1 0 89040 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_847
timestamp 1666464484
transform 1 0 96208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_851
timestamp 1666464484
transform 1 0 96656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_854
timestamp 1666464484
transform 1 0 96992 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_918
timestamp 1666464484
transform 1 0 104160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_922
timestamp 1666464484
transform 1 0 104608 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_925
timestamp 1666464484
transform 1 0 104944 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_989
timestamp 1666464484
transform 1 0 112112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_993
timestamp 1666464484
transform 1 0 112560 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_996
timestamp 1666464484
transform 1 0 112896 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1060
timestamp 1666464484
transform 1 0 120064 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1064
timestamp 1666464484
transform 1 0 120512 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1067
timestamp 1666464484
transform 1 0 120848 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1131
timestamp 1666464484
transform 1 0 128016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1135
timestamp 1666464484
transform 1 0 128464 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1138
timestamp 1666464484
transform 1 0 128800 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1202
timestamp 1666464484
transform 1 0 135968 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1206
timestamp 1666464484
transform 1 0 136416 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1209
timestamp 1666464484
transform 1 0 136752 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1273
timestamp 1666464484
transform 1 0 143920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1277
timestamp 1666464484
transform 1 0 144368 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1280
timestamp 1666464484
transform 1 0 144704 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1344
timestamp 1666464484
transform 1 0 151872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1348
timestamp 1666464484
transform 1 0 152320 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1351
timestamp 1666464484
transform 1 0 152656 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1415
timestamp 1666464484
transform 1 0 159824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1419
timestamp 1666464484
transform 1 0 160272 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1422
timestamp 1666464484
transform 1 0 160608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1486
timestamp 1666464484
transform 1 0 167776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1490
timestamp 1666464484
transform 1 0 168224 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1493
timestamp 1666464484
transform 1 0 168560 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1557
timestamp 1666464484
transform 1 0 175728 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1561
timestamp 1666464484
transform 1 0 176176 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_1564
timestamp 1666464484
transform 1 0 176512 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1580
timestamp 1666464484
transform 1 0 178304 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1666464484
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1666464484
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1666464484
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1666464484
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1666464484
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1666464484
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1666464484
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1666464484
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1666464484
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1666464484
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1666464484
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1666464484
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1666464484
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1666464484
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1666464484
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1666464484
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1666464484
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1666464484
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1666464484
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1666464484
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1666464484
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1666464484
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1666464484
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1666464484
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1666464484
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1666464484
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1666464484
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1666464484
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_676
timestamp 1666464484
transform 1 0 77056 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_740
timestamp 1666464484
transform 1 0 84224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_744
timestamp 1666464484
transform 1 0 84672 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_747
timestamp 1666464484
transform 1 0 85008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_811
timestamp 1666464484
transform 1 0 92176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_815
timestamp 1666464484
transform 1 0 92624 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_818
timestamp 1666464484
transform 1 0 92960 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_882
timestamp 1666464484
transform 1 0 100128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_886
timestamp 1666464484
transform 1 0 100576 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_889
timestamp 1666464484
transform 1 0 100912 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_953
timestamp 1666464484
transform 1 0 108080 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_957
timestamp 1666464484
transform 1 0 108528 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_960
timestamp 1666464484
transform 1 0 108864 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1024
timestamp 1666464484
transform 1 0 116032 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1028
timestamp 1666464484
transform 1 0 116480 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1031
timestamp 1666464484
transform 1 0 116816 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1095
timestamp 1666464484
transform 1 0 123984 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1099
timestamp 1666464484
transform 1 0 124432 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1102
timestamp 1666464484
transform 1 0 124768 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1166
timestamp 1666464484
transform 1 0 131936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1170
timestamp 1666464484
transform 1 0 132384 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1173
timestamp 1666464484
transform 1 0 132720 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1237
timestamp 1666464484
transform 1 0 139888 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1241
timestamp 1666464484
transform 1 0 140336 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1244
timestamp 1666464484
transform 1 0 140672 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1308
timestamp 1666464484
transform 1 0 147840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1312
timestamp 1666464484
transform 1 0 148288 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1315
timestamp 1666464484
transform 1 0 148624 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1379
timestamp 1666464484
transform 1 0 155792 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1383
timestamp 1666464484
transform 1 0 156240 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1386
timestamp 1666464484
transform 1 0 156576 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1450
timestamp 1666464484
transform 1 0 163744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1454
timestamp 1666464484
transform 1 0 164192 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1457
timestamp 1666464484
transform 1 0 164528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1521
timestamp 1666464484
transform 1 0 171696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1525
timestamp 1666464484
transform 1 0 172144 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_1528
timestamp 1666464484
transform 1 0 172480 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_1560
timestamp 1666464484
transform 1 0 176064 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1576
timestamp 1666464484
transform 1 0 177856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1580
timestamp 1666464484
transform 1 0 178304 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1666464484
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1666464484
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1666464484
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1666464484
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1666464484
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1666464484
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1666464484
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1666464484
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1666464484
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1666464484
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1666464484
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1666464484
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1666464484
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1666464484
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1666464484
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1666464484
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1666464484
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1666464484
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1666464484
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1666464484
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1666464484
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1666464484
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1666464484
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1666464484
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1666464484
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1666464484
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1666464484
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_641
timestamp 1666464484
transform 1 0 73136 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_705
timestamp 1666464484
transform 1 0 80304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_709
timestamp 1666464484
transform 1 0 80752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_712
timestamp 1666464484
transform 1 0 81088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_776
timestamp 1666464484
transform 1 0 88256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_780
timestamp 1666464484
transform 1 0 88704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_783
timestamp 1666464484
transform 1 0 89040 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_847
timestamp 1666464484
transform 1 0 96208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_851
timestamp 1666464484
transform 1 0 96656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_854
timestamp 1666464484
transform 1 0 96992 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_918
timestamp 1666464484
transform 1 0 104160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_922
timestamp 1666464484
transform 1 0 104608 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_925
timestamp 1666464484
transform 1 0 104944 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_989
timestamp 1666464484
transform 1 0 112112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_993
timestamp 1666464484
transform 1 0 112560 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_996
timestamp 1666464484
transform 1 0 112896 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1060
timestamp 1666464484
transform 1 0 120064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1064
timestamp 1666464484
transform 1 0 120512 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1067
timestamp 1666464484
transform 1 0 120848 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1131
timestamp 1666464484
transform 1 0 128016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1135
timestamp 1666464484
transform 1 0 128464 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1138
timestamp 1666464484
transform 1 0 128800 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1202
timestamp 1666464484
transform 1 0 135968 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1206
timestamp 1666464484
transform 1 0 136416 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1209
timestamp 1666464484
transform 1 0 136752 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1273
timestamp 1666464484
transform 1 0 143920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1277
timestamp 1666464484
transform 1 0 144368 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1280
timestamp 1666464484
transform 1 0 144704 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1344
timestamp 1666464484
transform 1 0 151872 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1348
timestamp 1666464484
transform 1 0 152320 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1351
timestamp 1666464484
transform 1 0 152656 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1415
timestamp 1666464484
transform 1 0 159824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1419
timestamp 1666464484
transform 1 0 160272 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1422
timestamp 1666464484
transform 1 0 160608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1486
timestamp 1666464484
transform 1 0 167776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1490
timestamp 1666464484
transform 1 0 168224 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1493
timestamp 1666464484
transform 1 0 168560 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1557
timestamp 1666464484
transform 1 0 175728 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1561
timestamp 1666464484
transform 1 0 176176 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_1564
timestamp 1666464484
transform 1 0 176512 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1580
timestamp 1666464484
transform 1 0 178304 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1666464484
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1666464484
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1666464484
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1666464484
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1666464484
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1666464484
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1666464484
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1666464484
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1666464484
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1666464484
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1666464484
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1666464484
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1666464484
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1666464484
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1666464484
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1666464484
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1666464484
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1666464484
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1666464484
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1666464484
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1666464484
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1666464484
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1666464484
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1666464484
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1666464484
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1666464484
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1666464484
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1666464484
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_676
timestamp 1666464484
transform 1 0 77056 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_740
timestamp 1666464484
transform 1 0 84224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_744
timestamp 1666464484
transform 1 0 84672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_747
timestamp 1666464484
transform 1 0 85008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_811
timestamp 1666464484
transform 1 0 92176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_815
timestamp 1666464484
transform 1 0 92624 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_818
timestamp 1666464484
transform 1 0 92960 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_882
timestamp 1666464484
transform 1 0 100128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_886
timestamp 1666464484
transform 1 0 100576 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_889
timestamp 1666464484
transform 1 0 100912 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_953
timestamp 1666464484
transform 1 0 108080 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_957
timestamp 1666464484
transform 1 0 108528 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_960
timestamp 1666464484
transform 1 0 108864 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1024
timestamp 1666464484
transform 1 0 116032 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1028
timestamp 1666464484
transform 1 0 116480 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1031
timestamp 1666464484
transform 1 0 116816 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1095
timestamp 1666464484
transform 1 0 123984 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1099
timestamp 1666464484
transform 1 0 124432 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1102
timestamp 1666464484
transform 1 0 124768 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1166
timestamp 1666464484
transform 1 0 131936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1170
timestamp 1666464484
transform 1 0 132384 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1173
timestamp 1666464484
transform 1 0 132720 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1237
timestamp 1666464484
transform 1 0 139888 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1241
timestamp 1666464484
transform 1 0 140336 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1244
timestamp 1666464484
transform 1 0 140672 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1308
timestamp 1666464484
transform 1 0 147840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1312
timestamp 1666464484
transform 1 0 148288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1315
timestamp 1666464484
transform 1 0 148624 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1379
timestamp 1666464484
transform 1 0 155792 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1383
timestamp 1666464484
transform 1 0 156240 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1386
timestamp 1666464484
transform 1 0 156576 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1450
timestamp 1666464484
transform 1 0 163744 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1454
timestamp 1666464484
transform 1 0 164192 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1457
timestamp 1666464484
transform 1 0 164528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1521
timestamp 1666464484
transform 1 0 171696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1525
timestamp 1666464484
transform 1 0 172144 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_1528
timestamp 1666464484
transform 1 0 172480 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_1560
timestamp 1666464484
transform 1 0 176064 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1576
timestamp 1666464484
transform 1 0 177856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1580
timestamp 1666464484
transform 1 0 178304 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1666464484
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1666464484
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1666464484
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1666464484
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1666464484
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1666464484
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1666464484
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1666464484
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1666464484
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1666464484
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1666464484
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1666464484
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1666464484
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1666464484
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1666464484
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1666464484
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1666464484
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1666464484
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1666464484
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1666464484
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1666464484
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1666464484
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1666464484
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1666464484
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1666464484
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1666464484
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1666464484
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_641
timestamp 1666464484
transform 1 0 73136 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_705
timestamp 1666464484
transform 1 0 80304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_709
timestamp 1666464484
transform 1 0 80752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_712
timestamp 1666464484
transform 1 0 81088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_776
timestamp 1666464484
transform 1 0 88256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_780
timestamp 1666464484
transform 1 0 88704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_783
timestamp 1666464484
transform 1 0 89040 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_847
timestamp 1666464484
transform 1 0 96208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_851
timestamp 1666464484
transform 1 0 96656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_854
timestamp 1666464484
transform 1 0 96992 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_918
timestamp 1666464484
transform 1 0 104160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_922
timestamp 1666464484
transform 1 0 104608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_925
timestamp 1666464484
transform 1 0 104944 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_989
timestamp 1666464484
transform 1 0 112112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_993
timestamp 1666464484
transform 1 0 112560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_996
timestamp 1666464484
transform 1 0 112896 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1060
timestamp 1666464484
transform 1 0 120064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1064
timestamp 1666464484
transform 1 0 120512 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1067
timestamp 1666464484
transform 1 0 120848 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1131
timestamp 1666464484
transform 1 0 128016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1135
timestamp 1666464484
transform 1 0 128464 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1138
timestamp 1666464484
transform 1 0 128800 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1202
timestamp 1666464484
transform 1 0 135968 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1206
timestamp 1666464484
transform 1 0 136416 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1209
timestamp 1666464484
transform 1 0 136752 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1273
timestamp 1666464484
transform 1 0 143920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1277
timestamp 1666464484
transform 1 0 144368 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1280
timestamp 1666464484
transform 1 0 144704 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1344
timestamp 1666464484
transform 1 0 151872 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1348
timestamp 1666464484
transform 1 0 152320 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1351
timestamp 1666464484
transform 1 0 152656 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1415
timestamp 1666464484
transform 1 0 159824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1419
timestamp 1666464484
transform 1 0 160272 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1422
timestamp 1666464484
transform 1 0 160608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1486
timestamp 1666464484
transform 1 0 167776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1490
timestamp 1666464484
transform 1 0 168224 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1493
timestamp 1666464484
transform 1 0 168560 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1557
timestamp 1666464484
transform 1 0 175728 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1561
timestamp 1666464484
transform 1 0 176176 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_1564
timestamp 1666464484
transform 1 0 176512 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1580
timestamp 1666464484
transform 1 0 178304 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1666464484
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1666464484
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1666464484
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1666464484
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1666464484
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1666464484
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1666464484
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1666464484
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1666464484
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1666464484
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1666464484
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1666464484
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1666464484
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1666464484
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1666464484
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1666464484
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1666464484
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1666464484
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1666464484
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1666464484
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1666464484
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1666464484
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1666464484
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1666464484
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1666464484
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1666464484
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1666464484
transform 1 0 76272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1666464484
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_676
timestamp 1666464484
transform 1 0 77056 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_740
timestamp 1666464484
transform 1 0 84224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_744
timestamp 1666464484
transform 1 0 84672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_747
timestamp 1666464484
transform 1 0 85008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_811
timestamp 1666464484
transform 1 0 92176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_815
timestamp 1666464484
transform 1 0 92624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_818
timestamp 1666464484
transform 1 0 92960 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_882
timestamp 1666464484
transform 1 0 100128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_886
timestamp 1666464484
transform 1 0 100576 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_889
timestamp 1666464484
transform 1 0 100912 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_953
timestamp 1666464484
transform 1 0 108080 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_957
timestamp 1666464484
transform 1 0 108528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_960
timestamp 1666464484
transform 1 0 108864 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1024
timestamp 1666464484
transform 1 0 116032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1028
timestamp 1666464484
transform 1 0 116480 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1031
timestamp 1666464484
transform 1 0 116816 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1095
timestamp 1666464484
transform 1 0 123984 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1099
timestamp 1666464484
transform 1 0 124432 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1102
timestamp 1666464484
transform 1 0 124768 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1166
timestamp 1666464484
transform 1 0 131936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1170
timestamp 1666464484
transform 1 0 132384 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1173
timestamp 1666464484
transform 1 0 132720 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1237
timestamp 1666464484
transform 1 0 139888 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1241
timestamp 1666464484
transform 1 0 140336 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1244
timestamp 1666464484
transform 1 0 140672 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1308
timestamp 1666464484
transform 1 0 147840 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1312
timestamp 1666464484
transform 1 0 148288 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1315
timestamp 1666464484
transform 1 0 148624 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1379
timestamp 1666464484
transform 1 0 155792 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1383
timestamp 1666464484
transform 1 0 156240 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1386
timestamp 1666464484
transform 1 0 156576 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1450
timestamp 1666464484
transform 1 0 163744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1454
timestamp 1666464484
transform 1 0 164192 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1457
timestamp 1666464484
transform 1 0 164528 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1521
timestamp 1666464484
transform 1 0 171696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1525
timestamp 1666464484
transform 1 0 172144 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_1528
timestamp 1666464484
transform 1 0 172480 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_1560
timestamp 1666464484
transform 1 0 176064 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1576
timestamp 1666464484
transform 1 0 177856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1580
timestamp 1666464484
transform 1 0 178304 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1666464484
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1666464484
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1666464484
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1666464484
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1666464484
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1666464484
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1666464484
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1666464484
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1666464484
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1666464484
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1666464484
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1666464484
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1666464484
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1666464484
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1666464484
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1666464484
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1666464484
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1666464484
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1666464484
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1666464484
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1666464484
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1666464484
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1666464484
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1666464484
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1666464484
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1666464484
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1666464484
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_641
timestamp 1666464484
transform 1 0 73136 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_705
timestamp 1666464484
transform 1 0 80304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_709
timestamp 1666464484
transform 1 0 80752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_712
timestamp 1666464484
transform 1 0 81088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_776
timestamp 1666464484
transform 1 0 88256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_780
timestamp 1666464484
transform 1 0 88704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_783
timestamp 1666464484
transform 1 0 89040 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_847
timestamp 1666464484
transform 1 0 96208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_851
timestamp 1666464484
transform 1 0 96656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_854
timestamp 1666464484
transform 1 0 96992 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_918
timestamp 1666464484
transform 1 0 104160 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_922
timestamp 1666464484
transform 1 0 104608 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_925
timestamp 1666464484
transform 1 0 104944 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_989
timestamp 1666464484
transform 1 0 112112 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_993
timestamp 1666464484
transform 1 0 112560 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_996
timestamp 1666464484
transform 1 0 112896 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1060
timestamp 1666464484
transform 1 0 120064 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1064
timestamp 1666464484
transform 1 0 120512 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1067
timestamp 1666464484
transform 1 0 120848 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1131
timestamp 1666464484
transform 1 0 128016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1135
timestamp 1666464484
transform 1 0 128464 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1138
timestamp 1666464484
transform 1 0 128800 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1202
timestamp 1666464484
transform 1 0 135968 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1206
timestamp 1666464484
transform 1 0 136416 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1209
timestamp 1666464484
transform 1 0 136752 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1273
timestamp 1666464484
transform 1 0 143920 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1277
timestamp 1666464484
transform 1 0 144368 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1280
timestamp 1666464484
transform 1 0 144704 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1344
timestamp 1666464484
transform 1 0 151872 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1348
timestamp 1666464484
transform 1 0 152320 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1351
timestamp 1666464484
transform 1 0 152656 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1415
timestamp 1666464484
transform 1 0 159824 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1419
timestamp 1666464484
transform 1 0 160272 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1422
timestamp 1666464484
transform 1 0 160608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1486
timestamp 1666464484
transform 1 0 167776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1490
timestamp 1666464484
transform 1 0 168224 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1493
timestamp 1666464484
transform 1 0 168560 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1557
timestamp 1666464484
transform 1 0 175728 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1561
timestamp 1666464484
transform 1 0 176176 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_1564
timestamp 1666464484
transform 1 0 176512 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1580
timestamp 1666464484
transform 1 0 178304 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1666464484
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1666464484
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1666464484
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1666464484
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1666464484
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1666464484
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1666464484
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1666464484
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1666464484
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1666464484
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1666464484
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1666464484
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1666464484
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1666464484
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1666464484
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1666464484
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1666464484
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1666464484
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1666464484
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1666464484
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1666464484
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1666464484
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1666464484
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1666464484
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1666464484
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1666464484
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1666464484
transform 1 0 76272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1666464484
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_676
timestamp 1666464484
transform 1 0 77056 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_740
timestamp 1666464484
transform 1 0 84224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_744
timestamp 1666464484
transform 1 0 84672 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_747
timestamp 1666464484
transform 1 0 85008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_811
timestamp 1666464484
transform 1 0 92176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_815
timestamp 1666464484
transform 1 0 92624 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_818
timestamp 1666464484
transform 1 0 92960 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_882
timestamp 1666464484
transform 1 0 100128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_886
timestamp 1666464484
transform 1 0 100576 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_889
timestamp 1666464484
transform 1 0 100912 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_953
timestamp 1666464484
transform 1 0 108080 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_957
timestamp 1666464484
transform 1 0 108528 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_960
timestamp 1666464484
transform 1 0 108864 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1024
timestamp 1666464484
transform 1 0 116032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1028
timestamp 1666464484
transform 1 0 116480 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1031
timestamp 1666464484
transform 1 0 116816 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1095
timestamp 1666464484
transform 1 0 123984 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1099
timestamp 1666464484
transform 1 0 124432 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1102
timestamp 1666464484
transform 1 0 124768 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1166
timestamp 1666464484
transform 1 0 131936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1170
timestamp 1666464484
transform 1 0 132384 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1173
timestamp 1666464484
transform 1 0 132720 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1237
timestamp 1666464484
transform 1 0 139888 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1241
timestamp 1666464484
transform 1 0 140336 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1244
timestamp 1666464484
transform 1 0 140672 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1308
timestamp 1666464484
transform 1 0 147840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1312
timestamp 1666464484
transform 1 0 148288 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1315
timestamp 1666464484
transform 1 0 148624 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1379
timestamp 1666464484
transform 1 0 155792 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1383
timestamp 1666464484
transform 1 0 156240 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1386
timestamp 1666464484
transform 1 0 156576 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1450
timestamp 1666464484
transform 1 0 163744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1454
timestamp 1666464484
transform 1 0 164192 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1457
timestamp 1666464484
transform 1 0 164528 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1521
timestamp 1666464484
transform 1 0 171696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1525
timestamp 1666464484
transform 1 0 172144 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_1528
timestamp 1666464484
transform 1 0 172480 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_1560
timestamp 1666464484
transform 1 0 176064 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1576
timestamp 1666464484
transform 1 0 177856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1580
timestamp 1666464484
transform 1 0 178304 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1666464484
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1666464484
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1666464484
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1666464484
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1666464484
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1666464484
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1666464484
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1666464484
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1666464484
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1666464484
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1666464484
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1666464484
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1666464484
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1666464484
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1666464484
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1666464484
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1666464484
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1666464484
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1666464484
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1666464484
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1666464484
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1666464484
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1666464484
transform 1 0 64400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1666464484
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1666464484
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1666464484
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1666464484
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_641
timestamp 1666464484
transform 1 0 73136 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_705
timestamp 1666464484
transform 1 0 80304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_709
timestamp 1666464484
transform 1 0 80752 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_712
timestamp 1666464484
transform 1 0 81088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_776
timestamp 1666464484
transform 1 0 88256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_780
timestamp 1666464484
transform 1 0 88704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_783
timestamp 1666464484
transform 1 0 89040 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_847
timestamp 1666464484
transform 1 0 96208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_851
timestamp 1666464484
transform 1 0 96656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_854
timestamp 1666464484
transform 1 0 96992 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_918
timestamp 1666464484
transform 1 0 104160 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_922
timestamp 1666464484
transform 1 0 104608 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_925
timestamp 1666464484
transform 1 0 104944 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_989
timestamp 1666464484
transform 1 0 112112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_993
timestamp 1666464484
transform 1 0 112560 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_996
timestamp 1666464484
transform 1 0 112896 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1060
timestamp 1666464484
transform 1 0 120064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1064
timestamp 1666464484
transform 1 0 120512 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1067
timestamp 1666464484
transform 1 0 120848 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1131
timestamp 1666464484
transform 1 0 128016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1135
timestamp 1666464484
transform 1 0 128464 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1138
timestamp 1666464484
transform 1 0 128800 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1202
timestamp 1666464484
transform 1 0 135968 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1206
timestamp 1666464484
transform 1 0 136416 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1209
timestamp 1666464484
transform 1 0 136752 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1273
timestamp 1666464484
transform 1 0 143920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1277
timestamp 1666464484
transform 1 0 144368 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1280
timestamp 1666464484
transform 1 0 144704 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1344
timestamp 1666464484
transform 1 0 151872 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1348
timestamp 1666464484
transform 1 0 152320 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1351
timestamp 1666464484
transform 1 0 152656 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1415
timestamp 1666464484
transform 1 0 159824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1419
timestamp 1666464484
transform 1 0 160272 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1422
timestamp 1666464484
transform 1 0 160608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1486
timestamp 1666464484
transform 1 0 167776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1490
timestamp 1666464484
transform 1 0 168224 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1493
timestamp 1666464484
transform 1 0 168560 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1557
timestamp 1666464484
transform 1 0 175728 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1561
timestamp 1666464484
transform 1 0 176176 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_1564
timestamp 1666464484
transform 1 0 176512 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1580
timestamp 1666464484
transform 1 0 178304 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1666464484
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1666464484
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1666464484
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1666464484
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1666464484
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1666464484
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1666464484
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1666464484
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1666464484
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1666464484
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1666464484
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1666464484
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1666464484
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1666464484
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1666464484
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1666464484
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1666464484
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1666464484
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1666464484
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1666464484
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1666464484
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1666464484
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1666464484
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1666464484
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1666464484
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1666464484
transform 1 0 69104 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_669
timestamp 1666464484
transform 1 0 76272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1666464484
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_676
timestamp 1666464484
transform 1 0 77056 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_740
timestamp 1666464484
transform 1 0 84224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_744
timestamp 1666464484
transform 1 0 84672 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_747
timestamp 1666464484
transform 1 0 85008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_811
timestamp 1666464484
transform 1 0 92176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_815
timestamp 1666464484
transform 1 0 92624 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_818
timestamp 1666464484
transform 1 0 92960 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_882
timestamp 1666464484
transform 1 0 100128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_886
timestamp 1666464484
transform 1 0 100576 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_889
timestamp 1666464484
transform 1 0 100912 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_953
timestamp 1666464484
transform 1 0 108080 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_957
timestamp 1666464484
transform 1 0 108528 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_960
timestamp 1666464484
transform 1 0 108864 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1024
timestamp 1666464484
transform 1 0 116032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1028
timestamp 1666464484
transform 1 0 116480 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1031
timestamp 1666464484
transform 1 0 116816 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1095
timestamp 1666464484
transform 1 0 123984 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1099
timestamp 1666464484
transform 1 0 124432 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1102
timestamp 1666464484
transform 1 0 124768 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1166
timestamp 1666464484
transform 1 0 131936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1170
timestamp 1666464484
transform 1 0 132384 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1173
timestamp 1666464484
transform 1 0 132720 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1237
timestamp 1666464484
transform 1 0 139888 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1241
timestamp 1666464484
transform 1 0 140336 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1244
timestamp 1666464484
transform 1 0 140672 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1308
timestamp 1666464484
transform 1 0 147840 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1312
timestamp 1666464484
transform 1 0 148288 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1315
timestamp 1666464484
transform 1 0 148624 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1379
timestamp 1666464484
transform 1 0 155792 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1383
timestamp 1666464484
transform 1 0 156240 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1386
timestamp 1666464484
transform 1 0 156576 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1450
timestamp 1666464484
transform 1 0 163744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1454
timestamp 1666464484
transform 1 0 164192 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1457
timestamp 1666464484
transform 1 0 164528 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1521
timestamp 1666464484
transform 1 0 171696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1525
timestamp 1666464484
transform 1 0 172144 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_1528
timestamp 1666464484
transform 1 0 172480 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1560
timestamp 1666464484
transform 1 0 176064 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1576
timestamp 1666464484
transform 1 0 177856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1580
timestamp 1666464484
transform 1 0 178304 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1666464484
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1666464484
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1666464484
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1666464484
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1666464484
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1666464484
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1666464484
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1666464484
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1666464484
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1666464484
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1666464484
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1666464484
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1666464484
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1666464484
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1666464484
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1666464484
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1666464484
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1666464484
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1666464484
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1666464484
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1666464484
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1666464484
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1666464484
transform 1 0 64400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1666464484
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1666464484
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1666464484
transform 1 0 72352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1666464484
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_641
timestamp 1666464484
transform 1 0 73136 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_705
timestamp 1666464484
transform 1 0 80304 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_709
timestamp 1666464484
transform 1 0 80752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_712
timestamp 1666464484
transform 1 0 81088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_776
timestamp 1666464484
transform 1 0 88256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_780
timestamp 1666464484
transform 1 0 88704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_783
timestamp 1666464484
transform 1 0 89040 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_847
timestamp 1666464484
transform 1 0 96208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_851
timestamp 1666464484
transform 1 0 96656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_854
timestamp 1666464484
transform 1 0 96992 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_918
timestamp 1666464484
transform 1 0 104160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_922
timestamp 1666464484
transform 1 0 104608 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_925
timestamp 1666464484
transform 1 0 104944 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_989
timestamp 1666464484
transform 1 0 112112 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_993
timestamp 1666464484
transform 1 0 112560 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_996
timestamp 1666464484
transform 1 0 112896 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1060
timestamp 1666464484
transform 1 0 120064 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1064
timestamp 1666464484
transform 1 0 120512 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1067
timestamp 1666464484
transform 1 0 120848 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1131
timestamp 1666464484
transform 1 0 128016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1135
timestamp 1666464484
transform 1 0 128464 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1138
timestamp 1666464484
transform 1 0 128800 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1202
timestamp 1666464484
transform 1 0 135968 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1206
timestamp 1666464484
transform 1 0 136416 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1209
timestamp 1666464484
transform 1 0 136752 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1273
timestamp 1666464484
transform 1 0 143920 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1277
timestamp 1666464484
transform 1 0 144368 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1280
timestamp 1666464484
transform 1 0 144704 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1344
timestamp 1666464484
transform 1 0 151872 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1348
timestamp 1666464484
transform 1 0 152320 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1351
timestamp 1666464484
transform 1 0 152656 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1415
timestamp 1666464484
transform 1 0 159824 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1419
timestamp 1666464484
transform 1 0 160272 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1422
timestamp 1666464484
transform 1 0 160608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1486
timestamp 1666464484
transform 1 0 167776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1490
timestamp 1666464484
transform 1 0 168224 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1493
timestamp 1666464484
transform 1 0 168560 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1557
timestamp 1666464484
transform 1 0 175728 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1561
timestamp 1666464484
transform 1 0 176176 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_1564
timestamp 1666464484
transform 1 0 176512 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1580
timestamp 1666464484
transform 1 0 178304 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1666464484
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1666464484
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1666464484
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1666464484
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1666464484
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1666464484
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1666464484
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1666464484
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1666464484
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1666464484
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1666464484
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1666464484
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1666464484
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1666464484
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1666464484
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1666464484
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1666464484
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1666464484
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1666464484
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1666464484
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1666464484
transform 1 0 53200 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1666464484
transform 1 0 60368 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1666464484
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1666464484
transform 1 0 68320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1666464484
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1666464484
transform 1 0 69104 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_669
timestamp 1666464484
transform 1 0 76272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1666464484
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_676
timestamp 1666464484
transform 1 0 77056 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_740
timestamp 1666464484
transform 1 0 84224 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_744
timestamp 1666464484
transform 1 0 84672 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_747
timestamp 1666464484
transform 1 0 85008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_811
timestamp 1666464484
transform 1 0 92176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_815
timestamp 1666464484
transform 1 0 92624 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_818
timestamp 1666464484
transform 1 0 92960 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_882
timestamp 1666464484
transform 1 0 100128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_886
timestamp 1666464484
transform 1 0 100576 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_889
timestamp 1666464484
transform 1 0 100912 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_953
timestamp 1666464484
transform 1 0 108080 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_957
timestamp 1666464484
transform 1 0 108528 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_960
timestamp 1666464484
transform 1 0 108864 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1024
timestamp 1666464484
transform 1 0 116032 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1028
timestamp 1666464484
transform 1 0 116480 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1031
timestamp 1666464484
transform 1 0 116816 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1095
timestamp 1666464484
transform 1 0 123984 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1099
timestamp 1666464484
transform 1 0 124432 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1102
timestamp 1666464484
transform 1 0 124768 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1166
timestamp 1666464484
transform 1 0 131936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1170
timestamp 1666464484
transform 1 0 132384 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1173
timestamp 1666464484
transform 1 0 132720 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1237
timestamp 1666464484
transform 1 0 139888 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1241
timestamp 1666464484
transform 1 0 140336 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1244
timestamp 1666464484
transform 1 0 140672 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1308
timestamp 1666464484
transform 1 0 147840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1312
timestamp 1666464484
transform 1 0 148288 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1315
timestamp 1666464484
transform 1 0 148624 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1379
timestamp 1666464484
transform 1 0 155792 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1383
timestamp 1666464484
transform 1 0 156240 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1386
timestamp 1666464484
transform 1 0 156576 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1450
timestamp 1666464484
transform 1 0 163744 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1454
timestamp 1666464484
transform 1 0 164192 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1457
timestamp 1666464484
transform 1 0 164528 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1521
timestamp 1666464484
transform 1 0 171696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1525
timestamp 1666464484
transform 1 0 172144 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_1528
timestamp 1666464484
transform 1 0 172480 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_1560
timestamp 1666464484
transform 1 0 176064 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1576
timestamp 1666464484
transform 1 0 177856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1580
timestamp 1666464484
transform 1 0 178304 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1666464484
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1666464484
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1666464484
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1666464484
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1666464484
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1666464484
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1666464484
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1666464484
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1666464484
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1666464484
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1666464484
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1666464484
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1666464484
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1666464484
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1666464484
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1666464484
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1666464484
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1666464484
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1666464484
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1666464484
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1666464484
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1666464484
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1666464484
transform 1 0 64400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1666464484
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1666464484
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1666464484
transform 1 0 72352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1666464484
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_641
timestamp 1666464484
transform 1 0 73136 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_705
timestamp 1666464484
transform 1 0 80304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_709
timestamp 1666464484
transform 1 0 80752 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_712
timestamp 1666464484
transform 1 0 81088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_776
timestamp 1666464484
transform 1 0 88256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_780
timestamp 1666464484
transform 1 0 88704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_783
timestamp 1666464484
transform 1 0 89040 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_847
timestamp 1666464484
transform 1 0 96208 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_851
timestamp 1666464484
transform 1 0 96656 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_854
timestamp 1666464484
transform 1 0 96992 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_918
timestamp 1666464484
transform 1 0 104160 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_922
timestamp 1666464484
transform 1 0 104608 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_925
timestamp 1666464484
transform 1 0 104944 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_989
timestamp 1666464484
transform 1 0 112112 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_993
timestamp 1666464484
transform 1 0 112560 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_996
timestamp 1666464484
transform 1 0 112896 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1060
timestamp 1666464484
transform 1 0 120064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1064
timestamp 1666464484
transform 1 0 120512 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1067
timestamp 1666464484
transform 1 0 120848 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1131
timestamp 1666464484
transform 1 0 128016 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1135
timestamp 1666464484
transform 1 0 128464 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1138
timestamp 1666464484
transform 1 0 128800 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1202
timestamp 1666464484
transform 1 0 135968 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1206
timestamp 1666464484
transform 1 0 136416 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1209
timestamp 1666464484
transform 1 0 136752 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1273
timestamp 1666464484
transform 1 0 143920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1277
timestamp 1666464484
transform 1 0 144368 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1280
timestamp 1666464484
transform 1 0 144704 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1344
timestamp 1666464484
transform 1 0 151872 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1348
timestamp 1666464484
transform 1 0 152320 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1351
timestamp 1666464484
transform 1 0 152656 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1415
timestamp 1666464484
transform 1 0 159824 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1419
timestamp 1666464484
transform 1 0 160272 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1422
timestamp 1666464484
transform 1 0 160608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1486
timestamp 1666464484
transform 1 0 167776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1490
timestamp 1666464484
transform 1 0 168224 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1493
timestamp 1666464484
transform 1 0 168560 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1557
timestamp 1666464484
transform 1 0 175728 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1561
timestamp 1666464484
transform 1 0 176176 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_1564
timestamp 1666464484
transform 1 0 176512 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1580
timestamp 1666464484
transform 1 0 178304 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1666464484
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1666464484
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1666464484
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1666464484
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1666464484
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1666464484
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1666464484
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1666464484
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1666464484
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1666464484
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1666464484
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1666464484
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1666464484
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1666464484
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1666464484
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1666464484
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1666464484
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1666464484
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_456
timestamp 1666464484
transform 1 0 52416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1666464484
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_463
timestamp 1666464484
transform 1 0 53200 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_527
timestamp 1666464484
transform 1 0 60368 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_531
timestamp 1666464484
transform 1 0 60816 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_534
timestamp 1666464484
transform 1 0 61152 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_598
timestamp 1666464484
transform 1 0 68320 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_602
timestamp 1666464484
transform 1 0 68768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_605
timestamp 1666464484
transform 1 0 69104 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_669
timestamp 1666464484
transform 1 0 76272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_673
timestamp 1666464484
transform 1 0 76720 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_676
timestamp 1666464484
transform 1 0 77056 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_740
timestamp 1666464484
transform 1 0 84224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_744
timestamp 1666464484
transform 1 0 84672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_747
timestamp 1666464484
transform 1 0 85008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_811
timestamp 1666464484
transform 1 0 92176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_815
timestamp 1666464484
transform 1 0 92624 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_818
timestamp 1666464484
transform 1 0 92960 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_882
timestamp 1666464484
transform 1 0 100128 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_886
timestamp 1666464484
transform 1 0 100576 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_889
timestamp 1666464484
transform 1 0 100912 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_953
timestamp 1666464484
transform 1 0 108080 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_957
timestamp 1666464484
transform 1 0 108528 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_960
timestamp 1666464484
transform 1 0 108864 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1024
timestamp 1666464484
transform 1 0 116032 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1028
timestamp 1666464484
transform 1 0 116480 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_1031
timestamp 1666464484
transform 1 0 116816 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1095
timestamp 1666464484
transform 1 0 123984 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1099
timestamp 1666464484
transform 1 0 124432 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_1102
timestamp 1666464484
transform 1 0 124768 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1166
timestamp 1666464484
transform 1 0 131936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1170
timestamp 1666464484
transform 1 0 132384 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_1173
timestamp 1666464484
transform 1 0 132720 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1237
timestamp 1666464484
transform 1 0 139888 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1241
timestamp 1666464484
transform 1 0 140336 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_1244
timestamp 1666464484
transform 1 0 140672 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1308
timestamp 1666464484
transform 1 0 147840 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1312
timestamp 1666464484
transform 1 0 148288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_1315
timestamp 1666464484
transform 1 0 148624 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1379
timestamp 1666464484
transform 1 0 155792 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1383
timestamp 1666464484
transform 1 0 156240 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_1386
timestamp 1666464484
transform 1 0 156576 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1450
timestamp 1666464484
transform 1 0 163744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1454
timestamp 1666464484
transform 1 0 164192 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_1457
timestamp 1666464484
transform 1 0 164528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1521
timestamp 1666464484
transform 1 0 171696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1525
timestamp 1666464484
transform 1 0 172144 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1528
timestamp 1666464484
transform 1 0 172480 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_1560
timestamp 1666464484
transform 1 0 176064 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1576
timestamp 1666464484
transform 1 0 177856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1580
timestamp 1666464484
transform 1 0 178304 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1666464484
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1666464484
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1666464484
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1666464484
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1666464484
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1666464484
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1666464484
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1666464484
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1666464484
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1666464484
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1666464484
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1666464484
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1666464484
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1666464484
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1666464484
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1666464484
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1666464484
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1666464484
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_428
timestamp 1666464484
transform 1 0 49280 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_492
timestamp 1666464484
transform 1 0 56448 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1666464484
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_499
timestamp 1666464484
transform 1 0 57232 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_563
timestamp 1666464484
transform 1 0 64400 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_567
timestamp 1666464484
transform 1 0 64848 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_570
timestamp 1666464484
transform 1 0 65184 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_634
timestamp 1666464484
transform 1 0 72352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_638
timestamp 1666464484
transform 1 0 72800 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_641
timestamp 1666464484
transform 1 0 73136 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_705
timestamp 1666464484
transform 1 0 80304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_709
timestamp 1666464484
transform 1 0 80752 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_712
timestamp 1666464484
transform 1 0 81088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_776
timestamp 1666464484
transform 1 0 88256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_780
timestamp 1666464484
transform 1 0 88704 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_783
timestamp 1666464484
transform 1 0 89040 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_847
timestamp 1666464484
transform 1 0 96208 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_851
timestamp 1666464484
transform 1 0 96656 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_854
timestamp 1666464484
transform 1 0 96992 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_918
timestamp 1666464484
transform 1 0 104160 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_922
timestamp 1666464484
transform 1 0 104608 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_925
timestamp 1666464484
transform 1 0 104944 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_989
timestamp 1666464484
transform 1 0 112112 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_993
timestamp 1666464484
transform 1 0 112560 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_996
timestamp 1666464484
transform 1 0 112896 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_1060
timestamp 1666464484
transform 1 0 120064 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1064
timestamp 1666464484
transform 1 0 120512 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_1067
timestamp 1666464484
transform 1 0 120848 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_1131
timestamp 1666464484
transform 1 0 128016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1135
timestamp 1666464484
transform 1 0 128464 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_1138
timestamp 1666464484
transform 1 0 128800 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_1202
timestamp 1666464484
transform 1 0 135968 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1206
timestamp 1666464484
transform 1 0 136416 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_1209
timestamp 1666464484
transform 1 0 136752 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_1273
timestamp 1666464484
transform 1 0 143920 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1277
timestamp 1666464484
transform 1 0 144368 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_1280
timestamp 1666464484
transform 1 0 144704 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_1344
timestamp 1666464484
transform 1 0 151872 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1348
timestamp 1666464484
transform 1 0 152320 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_1351
timestamp 1666464484
transform 1 0 152656 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_1415
timestamp 1666464484
transform 1 0 159824 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1419
timestamp 1666464484
transform 1 0 160272 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_1422
timestamp 1666464484
transform 1 0 160608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_1486
timestamp 1666464484
transform 1 0 167776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1490
timestamp 1666464484
transform 1 0 168224 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_1493
timestamp 1666464484
transform 1 0 168560 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_1557
timestamp 1666464484
transform 1 0 175728 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1561
timestamp 1666464484
transform 1 0 176176 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_1564
timestamp 1666464484
transform 1 0 176512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1580
timestamp 1666464484
transform 1 0 178304 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1666464484
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1666464484
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1666464484
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1666464484
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1666464484
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1666464484
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1666464484
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1666464484
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1666464484
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1666464484
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1666464484
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1666464484
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1666464484
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1666464484
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1666464484
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1666464484
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1666464484
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1666464484
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1666464484
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1666464484
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_463
timestamp 1666464484
transform 1 0 53200 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_527
timestamp 1666464484
transform 1 0 60368 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 60816 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_534
timestamp 1666464484
transform 1 0 61152 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_598
timestamp 1666464484
transform 1 0 68320 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_602
timestamp 1666464484
transform 1 0 68768 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_605
timestamp 1666464484
transform 1 0 69104 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_669
timestamp 1666464484
transform 1 0 76272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_673
timestamp 1666464484
transform 1 0 76720 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_676
timestamp 1666464484
transform 1 0 77056 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_740
timestamp 1666464484
transform 1 0 84224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_744
timestamp 1666464484
transform 1 0 84672 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_747
timestamp 1666464484
transform 1 0 85008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_811
timestamp 1666464484
transform 1 0 92176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_815
timestamp 1666464484
transform 1 0 92624 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_818
timestamp 1666464484
transform 1 0 92960 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_882
timestamp 1666464484
transform 1 0 100128 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_886
timestamp 1666464484
transform 1 0 100576 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_889
timestamp 1666464484
transform 1 0 100912 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_953
timestamp 1666464484
transform 1 0 108080 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_957
timestamp 1666464484
transform 1 0 108528 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_960
timestamp 1666464484
transform 1 0 108864 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1024
timestamp 1666464484
transform 1 0 116032 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1028
timestamp 1666464484
transform 1 0 116480 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_1031
timestamp 1666464484
transform 1 0 116816 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1095
timestamp 1666464484
transform 1 0 123984 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1099
timestamp 1666464484
transform 1 0 124432 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_1102
timestamp 1666464484
transform 1 0 124768 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1166
timestamp 1666464484
transform 1 0 131936 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1170
timestamp 1666464484
transform 1 0 132384 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_1173
timestamp 1666464484
transform 1 0 132720 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1237
timestamp 1666464484
transform 1 0 139888 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1241
timestamp 1666464484
transform 1 0 140336 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_1244
timestamp 1666464484
transform 1 0 140672 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1308
timestamp 1666464484
transform 1 0 147840 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1312
timestamp 1666464484
transform 1 0 148288 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_1315
timestamp 1666464484
transform 1 0 148624 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1379
timestamp 1666464484
transform 1 0 155792 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1383
timestamp 1666464484
transform 1 0 156240 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_1386
timestamp 1666464484
transform 1 0 156576 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1450
timestamp 1666464484
transform 1 0 163744 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1454
timestamp 1666464484
transform 1 0 164192 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_1457
timestamp 1666464484
transform 1 0 164528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1521
timestamp 1666464484
transform 1 0 171696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1525
timestamp 1666464484
transform 1 0 172144 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_1528
timestamp 1666464484
transform 1 0 172480 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_1560
timestamp 1666464484
transform 1 0 176064 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1576
timestamp 1666464484
transform 1 0 177856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1580
timestamp 1666464484
transform 1 0 178304 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1666464484
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1666464484
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1666464484
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1666464484
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1666464484
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1666464484
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1666464484
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1666464484
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1666464484
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1666464484
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1666464484
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1666464484
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1666464484
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1666464484
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1666464484
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1666464484
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1666464484
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1666464484
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_428
timestamp 1666464484
transform 1 0 49280 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_492
timestamp 1666464484
transform 1 0 56448 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1666464484
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_499
timestamp 1666464484
transform 1 0 57232 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_563
timestamp 1666464484
transform 1 0 64400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_567
timestamp 1666464484
transform 1 0 64848 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_570
timestamp 1666464484
transform 1 0 65184 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_634
timestamp 1666464484
transform 1 0 72352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_638
timestamp 1666464484
transform 1 0 72800 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_641
timestamp 1666464484
transform 1 0 73136 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_705
timestamp 1666464484
transform 1 0 80304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_709
timestamp 1666464484
transform 1 0 80752 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_712
timestamp 1666464484
transform 1 0 81088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_776
timestamp 1666464484
transform 1 0 88256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_780
timestamp 1666464484
transform 1 0 88704 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_783
timestamp 1666464484
transform 1 0 89040 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_847
timestamp 1666464484
transform 1 0 96208 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_851
timestamp 1666464484
transform 1 0 96656 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_854
timestamp 1666464484
transform 1 0 96992 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_918
timestamp 1666464484
transform 1 0 104160 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_922
timestamp 1666464484
transform 1 0 104608 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_925
timestamp 1666464484
transform 1 0 104944 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_989
timestamp 1666464484
transform 1 0 112112 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_993
timestamp 1666464484
transform 1 0 112560 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_996
timestamp 1666464484
transform 1 0 112896 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1060
timestamp 1666464484
transform 1 0 120064 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1064
timestamp 1666464484
transform 1 0 120512 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_1067
timestamp 1666464484
transform 1 0 120848 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1131
timestamp 1666464484
transform 1 0 128016 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1135
timestamp 1666464484
transform 1 0 128464 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_1138
timestamp 1666464484
transform 1 0 128800 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1202
timestamp 1666464484
transform 1 0 135968 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1206
timestamp 1666464484
transform 1 0 136416 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_1209
timestamp 1666464484
transform 1 0 136752 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1273
timestamp 1666464484
transform 1 0 143920 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1277
timestamp 1666464484
transform 1 0 144368 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_1280
timestamp 1666464484
transform 1 0 144704 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1344
timestamp 1666464484
transform 1 0 151872 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1348
timestamp 1666464484
transform 1 0 152320 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_1351
timestamp 1666464484
transform 1 0 152656 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1415
timestamp 1666464484
transform 1 0 159824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1419
timestamp 1666464484
transform 1 0 160272 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_1422
timestamp 1666464484
transform 1 0 160608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1486
timestamp 1666464484
transform 1 0 167776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1490
timestamp 1666464484
transform 1 0 168224 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_1493
timestamp 1666464484
transform 1 0 168560 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1557
timestamp 1666464484
transform 1 0 175728 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1561
timestamp 1666464484
transform 1 0 176176 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_1564
timestamp 1666464484
transform 1 0 176512 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1580
timestamp 1666464484
transform 1 0 178304 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1666464484
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1666464484
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1666464484
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1666464484
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1666464484
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1666464484
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1666464484
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1666464484
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1666464484
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1666464484
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1666464484
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1666464484
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1666464484
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1666464484
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1666464484
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1666464484
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1666464484
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_392
timestamp 1666464484
transform 1 0 45248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_456
timestamp 1666464484
transform 1 0 52416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1666464484
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_463
timestamp 1666464484
transform 1 0 53200 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_527
timestamp 1666464484
transform 1 0 60368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_531
timestamp 1666464484
transform 1 0 60816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_534
timestamp 1666464484
transform 1 0 61152 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_598
timestamp 1666464484
transform 1 0 68320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_602
timestamp 1666464484
transform 1 0 68768 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_605
timestamp 1666464484
transform 1 0 69104 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_669
timestamp 1666464484
transform 1 0 76272 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_673
timestamp 1666464484
transform 1 0 76720 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_676
timestamp 1666464484
transform 1 0 77056 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_740
timestamp 1666464484
transform 1 0 84224 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_744
timestamp 1666464484
transform 1 0 84672 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_747
timestamp 1666464484
transform 1 0 85008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_811
timestamp 1666464484
transform 1 0 92176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_815
timestamp 1666464484
transform 1 0 92624 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_818
timestamp 1666464484
transform 1 0 92960 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_882
timestamp 1666464484
transform 1 0 100128 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_886
timestamp 1666464484
transform 1 0 100576 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_889
timestamp 1666464484
transform 1 0 100912 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_953
timestamp 1666464484
transform 1 0 108080 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_957
timestamp 1666464484
transform 1 0 108528 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_960
timestamp 1666464484
transform 1 0 108864 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1024
timestamp 1666464484
transform 1 0 116032 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1028
timestamp 1666464484
transform 1 0 116480 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_1031
timestamp 1666464484
transform 1 0 116816 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1095
timestamp 1666464484
transform 1 0 123984 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1099
timestamp 1666464484
transform 1 0 124432 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_1102
timestamp 1666464484
transform 1 0 124768 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1166
timestamp 1666464484
transform 1 0 131936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1170
timestamp 1666464484
transform 1 0 132384 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_1173
timestamp 1666464484
transform 1 0 132720 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1237
timestamp 1666464484
transform 1 0 139888 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1241
timestamp 1666464484
transform 1 0 140336 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_1244
timestamp 1666464484
transform 1 0 140672 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1308
timestamp 1666464484
transform 1 0 147840 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1312
timestamp 1666464484
transform 1 0 148288 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_1315
timestamp 1666464484
transform 1 0 148624 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1379
timestamp 1666464484
transform 1 0 155792 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1383
timestamp 1666464484
transform 1 0 156240 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_1386
timestamp 1666464484
transform 1 0 156576 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1450
timestamp 1666464484
transform 1 0 163744 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1454
timestamp 1666464484
transform 1 0 164192 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_1457
timestamp 1666464484
transform 1 0 164528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1521
timestamp 1666464484
transform 1 0 171696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1525
timestamp 1666464484
transform 1 0 172144 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_1528
timestamp 1666464484
transform 1 0 172480 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_1560
timestamp 1666464484
transform 1 0 176064 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1576
timestamp 1666464484
transform 1 0 177856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1580
timestamp 1666464484
transform 1 0 178304 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1666464484
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1666464484
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1666464484
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1666464484
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1666464484
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1666464484
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1666464484
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1666464484
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1666464484
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1666464484
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1666464484
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1666464484
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1666464484
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1666464484
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1666464484
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_357
timestamp 1666464484
transform 1 0 41328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_421
timestamp 1666464484
transform 1 0 48496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_425
timestamp 1666464484
transform 1 0 48944 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1666464484
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1666464484
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1666464484
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_499
timestamp 1666464484
transform 1 0 57232 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_563
timestamp 1666464484
transform 1 0 64400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_567
timestamp 1666464484
transform 1 0 64848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_570
timestamp 1666464484
transform 1 0 65184 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_634
timestamp 1666464484
transform 1 0 72352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_638
timestamp 1666464484
transform 1 0 72800 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_641
timestamp 1666464484
transform 1 0 73136 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_705
timestamp 1666464484
transform 1 0 80304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_709
timestamp 1666464484
transform 1 0 80752 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_712
timestamp 1666464484
transform 1 0 81088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_776
timestamp 1666464484
transform 1 0 88256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_780
timestamp 1666464484
transform 1 0 88704 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_783
timestamp 1666464484
transform 1 0 89040 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_847
timestamp 1666464484
transform 1 0 96208 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_851
timestamp 1666464484
transform 1 0 96656 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_854
timestamp 1666464484
transform 1 0 96992 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_918
timestamp 1666464484
transform 1 0 104160 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_922
timestamp 1666464484
transform 1 0 104608 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_925
timestamp 1666464484
transform 1 0 104944 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_989
timestamp 1666464484
transform 1 0 112112 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_993
timestamp 1666464484
transform 1 0 112560 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_996
timestamp 1666464484
transform 1 0 112896 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1060
timestamp 1666464484
transform 1 0 120064 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1064
timestamp 1666464484
transform 1 0 120512 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_1067
timestamp 1666464484
transform 1 0 120848 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1131
timestamp 1666464484
transform 1 0 128016 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1135
timestamp 1666464484
transform 1 0 128464 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_1138
timestamp 1666464484
transform 1 0 128800 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1202
timestamp 1666464484
transform 1 0 135968 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1206
timestamp 1666464484
transform 1 0 136416 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_1209
timestamp 1666464484
transform 1 0 136752 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1273
timestamp 1666464484
transform 1 0 143920 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1277
timestamp 1666464484
transform 1 0 144368 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_1280
timestamp 1666464484
transform 1 0 144704 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1344
timestamp 1666464484
transform 1 0 151872 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1348
timestamp 1666464484
transform 1 0 152320 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_1351
timestamp 1666464484
transform 1 0 152656 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1415
timestamp 1666464484
transform 1 0 159824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1419
timestamp 1666464484
transform 1 0 160272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_1422
timestamp 1666464484
transform 1 0 160608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1486
timestamp 1666464484
transform 1 0 167776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1490
timestamp 1666464484
transform 1 0 168224 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_1493
timestamp 1666464484
transform 1 0 168560 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_1557
timestamp 1666464484
transform 1 0 175728 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1561
timestamp 1666464484
transform 1 0 176176 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_1564
timestamp 1666464484
transform 1 0 176512 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1580
timestamp 1666464484
transform 1 0 178304 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_2
timestamp 1666464484
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1666464484
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1666464484
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1666464484
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1666464484
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1666464484
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1666464484
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1666464484
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1666464484
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1666464484
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1666464484
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1666464484
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1666464484
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1666464484
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1666464484
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1666464484
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1666464484
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1666464484
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_456
timestamp 1666464484
transform 1 0 52416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1666464484
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_463
timestamp 1666464484
transform 1 0 53200 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_527
timestamp 1666464484
transform 1 0 60368 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 60816 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_534
timestamp 1666464484
transform 1 0 61152 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_598
timestamp 1666464484
transform 1 0 68320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_602
timestamp 1666464484
transform 1 0 68768 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_605
timestamp 1666464484
transform 1 0 69104 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_669
timestamp 1666464484
transform 1 0 76272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_673
timestamp 1666464484
transform 1 0 76720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_676
timestamp 1666464484
transform 1 0 77056 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_740
timestamp 1666464484
transform 1 0 84224 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_744
timestamp 1666464484
transform 1 0 84672 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_747
timestamp 1666464484
transform 1 0 85008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_811
timestamp 1666464484
transform 1 0 92176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_815
timestamp 1666464484
transform 1 0 92624 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_818
timestamp 1666464484
transform 1 0 92960 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_882
timestamp 1666464484
transform 1 0 100128 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_886
timestamp 1666464484
transform 1 0 100576 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_889
timestamp 1666464484
transform 1 0 100912 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_953
timestamp 1666464484
transform 1 0 108080 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_957
timestamp 1666464484
transform 1 0 108528 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_960
timestamp 1666464484
transform 1 0 108864 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1024
timestamp 1666464484
transform 1 0 116032 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1028
timestamp 1666464484
transform 1 0 116480 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_1031
timestamp 1666464484
transform 1 0 116816 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1095
timestamp 1666464484
transform 1 0 123984 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1099
timestamp 1666464484
transform 1 0 124432 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_1102
timestamp 1666464484
transform 1 0 124768 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1166
timestamp 1666464484
transform 1 0 131936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1170
timestamp 1666464484
transform 1 0 132384 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_1173
timestamp 1666464484
transform 1 0 132720 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1237
timestamp 1666464484
transform 1 0 139888 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1241
timestamp 1666464484
transform 1 0 140336 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_1244
timestamp 1666464484
transform 1 0 140672 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1308
timestamp 1666464484
transform 1 0 147840 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1312
timestamp 1666464484
transform 1 0 148288 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_1315
timestamp 1666464484
transform 1 0 148624 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1379
timestamp 1666464484
transform 1 0 155792 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1383
timestamp 1666464484
transform 1 0 156240 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_1386
timestamp 1666464484
transform 1 0 156576 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1450
timestamp 1666464484
transform 1 0 163744 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1454
timestamp 1666464484
transform 1 0 164192 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_1457
timestamp 1666464484
transform 1 0 164528 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1521
timestamp 1666464484
transform 1 0 171696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1525
timestamp 1666464484
transform 1 0 172144 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_1528
timestamp 1666464484
transform 1 0 172480 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_1560
timestamp 1666464484
transform 1 0 176064 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1576
timestamp 1666464484
transform 1 0 177856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1580
timestamp 1666464484
transform 1 0 178304 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1666464484
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1666464484
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1666464484
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1666464484
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1666464484
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1666464484
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1666464484
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1666464484
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1666464484
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1666464484
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1666464484
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1666464484
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1666464484
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1666464484
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1666464484
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_357
timestamp 1666464484
transform 1 0 41328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_421
timestamp 1666464484
transform 1 0 48496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1666464484
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1666464484
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_492
timestamp 1666464484
transform 1 0 56448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1666464484
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_499
timestamp 1666464484
transform 1 0 57232 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_563
timestamp 1666464484
transform 1 0 64400 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_567
timestamp 1666464484
transform 1 0 64848 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_570
timestamp 1666464484
transform 1 0 65184 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_634
timestamp 1666464484
transform 1 0 72352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_638
timestamp 1666464484
transform 1 0 72800 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_641
timestamp 1666464484
transform 1 0 73136 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_705
timestamp 1666464484
transform 1 0 80304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_709
timestamp 1666464484
transform 1 0 80752 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_712
timestamp 1666464484
transform 1 0 81088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_776
timestamp 1666464484
transform 1 0 88256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_780
timestamp 1666464484
transform 1 0 88704 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_783
timestamp 1666464484
transform 1 0 89040 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_847
timestamp 1666464484
transform 1 0 96208 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_851
timestamp 1666464484
transform 1 0 96656 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_854
timestamp 1666464484
transform 1 0 96992 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_918
timestamp 1666464484
transform 1 0 104160 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_922
timestamp 1666464484
transform 1 0 104608 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_925
timestamp 1666464484
transform 1 0 104944 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_989
timestamp 1666464484
transform 1 0 112112 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_993
timestamp 1666464484
transform 1 0 112560 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_996
timestamp 1666464484
transform 1 0 112896 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1060
timestamp 1666464484
transform 1 0 120064 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1064
timestamp 1666464484
transform 1 0 120512 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_1067
timestamp 1666464484
transform 1 0 120848 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1131
timestamp 1666464484
transform 1 0 128016 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1135
timestamp 1666464484
transform 1 0 128464 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_1138
timestamp 1666464484
transform 1 0 128800 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1202
timestamp 1666464484
transform 1 0 135968 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1206
timestamp 1666464484
transform 1 0 136416 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_1209
timestamp 1666464484
transform 1 0 136752 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1273
timestamp 1666464484
transform 1 0 143920 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1277
timestamp 1666464484
transform 1 0 144368 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_1280
timestamp 1666464484
transform 1 0 144704 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1344
timestamp 1666464484
transform 1 0 151872 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1348
timestamp 1666464484
transform 1 0 152320 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_1351
timestamp 1666464484
transform 1 0 152656 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1415
timestamp 1666464484
transform 1 0 159824 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1419
timestamp 1666464484
transform 1 0 160272 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_1422
timestamp 1666464484
transform 1 0 160608 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1486
timestamp 1666464484
transform 1 0 167776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1490
timestamp 1666464484
transform 1 0 168224 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_1493
timestamp 1666464484
transform 1 0 168560 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_1557
timestamp 1666464484
transform 1 0 175728 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1561
timestamp 1666464484
transform 1 0 176176 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_1564
timestamp 1666464484
transform 1 0 176512 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1580
timestamp 1666464484
transform 1 0 178304 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1666464484
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1666464484
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1666464484
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1666464484
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1666464484
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1666464484
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1666464484
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1666464484
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1666464484
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1666464484
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1666464484
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1666464484
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1666464484
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1666464484
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1666464484
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1666464484
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1666464484
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_392
timestamp 1666464484
transform 1 0 45248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_456
timestamp 1666464484
transform 1 0 52416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1666464484
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_463
timestamp 1666464484
transform 1 0 53200 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_527
timestamp 1666464484
transform 1 0 60368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 60816 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_534
timestamp 1666464484
transform 1 0 61152 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_598
timestamp 1666464484
transform 1 0 68320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_602
timestamp 1666464484
transform 1 0 68768 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_605
timestamp 1666464484
transform 1 0 69104 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_669
timestamp 1666464484
transform 1 0 76272 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_673
timestamp 1666464484
transform 1 0 76720 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_676
timestamp 1666464484
transform 1 0 77056 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_740
timestamp 1666464484
transform 1 0 84224 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_744
timestamp 1666464484
transform 1 0 84672 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_747
timestamp 1666464484
transform 1 0 85008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_811
timestamp 1666464484
transform 1 0 92176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_815
timestamp 1666464484
transform 1 0 92624 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_818
timestamp 1666464484
transform 1 0 92960 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_882
timestamp 1666464484
transform 1 0 100128 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_886
timestamp 1666464484
transform 1 0 100576 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_889
timestamp 1666464484
transform 1 0 100912 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_953
timestamp 1666464484
transform 1 0 108080 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_957
timestamp 1666464484
transform 1 0 108528 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_960
timestamp 1666464484
transform 1 0 108864 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1024
timestamp 1666464484
transform 1 0 116032 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1028
timestamp 1666464484
transform 1 0 116480 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_1031
timestamp 1666464484
transform 1 0 116816 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1095
timestamp 1666464484
transform 1 0 123984 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1099
timestamp 1666464484
transform 1 0 124432 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_1102
timestamp 1666464484
transform 1 0 124768 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1166
timestamp 1666464484
transform 1 0 131936 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1170
timestamp 1666464484
transform 1 0 132384 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_1173
timestamp 1666464484
transform 1 0 132720 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1237
timestamp 1666464484
transform 1 0 139888 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1241
timestamp 1666464484
transform 1 0 140336 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_1244
timestamp 1666464484
transform 1 0 140672 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1308
timestamp 1666464484
transform 1 0 147840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1312
timestamp 1666464484
transform 1 0 148288 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_1315
timestamp 1666464484
transform 1 0 148624 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1379
timestamp 1666464484
transform 1 0 155792 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1383
timestamp 1666464484
transform 1 0 156240 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_1386
timestamp 1666464484
transform 1 0 156576 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1450
timestamp 1666464484
transform 1 0 163744 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1454
timestamp 1666464484
transform 1 0 164192 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_1457
timestamp 1666464484
transform 1 0 164528 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1521
timestamp 1666464484
transform 1 0 171696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1525
timestamp 1666464484
transform 1 0 172144 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_1528
timestamp 1666464484
transform 1 0 172480 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_1560
timestamp 1666464484
transform 1 0 176064 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1576
timestamp 1666464484
transform 1 0 177856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1580
timestamp 1666464484
transform 1 0 178304 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1666464484
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1666464484
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1666464484
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1666464484
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1666464484
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1666464484
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1666464484
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1666464484
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1666464484
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1666464484
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1666464484
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1666464484
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1666464484
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1666464484
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1666464484
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_357
timestamp 1666464484
transform 1 0 41328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_421
timestamp 1666464484
transform 1 0 48496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1666464484
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1666464484
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1666464484
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1666464484
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_499
timestamp 1666464484
transform 1 0 57232 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_563
timestamp 1666464484
transform 1 0 64400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_567
timestamp 1666464484
transform 1 0 64848 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_570
timestamp 1666464484
transform 1 0 65184 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_634
timestamp 1666464484
transform 1 0 72352 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_638
timestamp 1666464484
transform 1 0 72800 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_641
timestamp 1666464484
transform 1 0 73136 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_705
timestamp 1666464484
transform 1 0 80304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_709
timestamp 1666464484
transform 1 0 80752 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_712
timestamp 1666464484
transform 1 0 81088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_776
timestamp 1666464484
transform 1 0 88256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_780
timestamp 1666464484
transform 1 0 88704 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_783
timestamp 1666464484
transform 1 0 89040 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_847
timestamp 1666464484
transform 1 0 96208 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_851
timestamp 1666464484
transform 1 0 96656 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_854
timestamp 1666464484
transform 1 0 96992 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_918
timestamp 1666464484
transform 1 0 104160 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_922
timestamp 1666464484
transform 1 0 104608 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_925
timestamp 1666464484
transform 1 0 104944 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_989
timestamp 1666464484
transform 1 0 112112 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_993
timestamp 1666464484
transform 1 0 112560 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_996
timestamp 1666464484
transform 1 0 112896 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1060
timestamp 1666464484
transform 1 0 120064 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1064
timestamp 1666464484
transform 1 0 120512 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_1067
timestamp 1666464484
transform 1 0 120848 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1131
timestamp 1666464484
transform 1 0 128016 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1135
timestamp 1666464484
transform 1 0 128464 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_1138
timestamp 1666464484
transform 1 0 128800 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1202
timestamp 1666464484
transform 1 0 135968 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1206
timestamp 1666464484
transform 1 0 136416 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_1209
timestamp 1666464484
transform 1 0 136752 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1273
timestamp 1666464484
transform 1 0 143920 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1277
timestamp 1666464484
transform 1 0 144368 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_1280
timestamp 1666464484
transform 1 0 144704 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1344
timestamp 1666464484
transform 1 0 151872 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1348
timestamp 1666464484
transform 1 0 152320 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_1351
timestamp 1666464484
transform 1 0 152656 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1415
timestamp 1666464484
transform 1 0 159824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1419
timestamp 1666464484
transform 1 0 160272 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_1422
timestamp 1666464484
transform 1 0 160608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1486
timestamp 1666464484
transform 1 0 167776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1490
timestamp 1666464484
transform 1 0 168224 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_1493
timestamp 1666464484
transform 1 0 168560 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_1557
timestamp 1666464484
transform 1 0 175728 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1561
timestamp 1666464484
transform 1 0 176176 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_1564
timestamp 1666464484
transform 1 0 176512 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1580
timestamp 1666464484
transform 1 0 178304 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1666464484
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1666464484
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1666464484
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1666464484
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1666464484
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1666464484
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1666464484
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1666464484
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1666464484
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1666464484
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1666464484
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1666464484
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1666464484
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1666464484
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1666464484
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1666464484
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1666464484
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_392
timestamp 1666464484
transform 1 0 45248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_456
timestamp 1666464484
transform 1 0 52416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1666464484
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_463
timestamp 1666464484
transform 1 0 53200 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_527
timestamp 1666464484
transform 1 0 60368 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 60816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_534
timestamp 1666464484
transform 1 0 61152 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_598
timestamp 1666464484
transform 1 0 68320 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_602
timestamp 1666464484
transform 1 0 68768 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_605
timestamp 1666464484
transform 1 0 69104 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_669
timestamp 1666464484
transform 1 0 76272 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_673
timestamp 1666464484
transform 1 0 76720 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_676
timestamp 1666464484
transform 1 0 77056 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_740
timestamp 1666464484
transform 1 0 84224 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_744
timestamp 1666464484
transform 1 0 84672 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_747
timestamp 1666464484
transform 1 0 85008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_811
timestamp 1666464484
transform 1 0 92176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_815
timestamp 1666464484
transform 1 0 92624 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_818
timestamp 1666464484
transform 1 0 92960 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_882
timestamp 1666464484
transform 1 0 100128 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_886
timestamp 1666464484
transform 1 0 100576 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_889
timestamp 1666464484
transform 1 0 100912 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_953
timestamp 1666464484
transform 1 0 108080 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_957
timestamp 1666464484
transform 1 0 108528 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_960
timestamp 1666464484
transform 1 0 108864 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1024
timestamp 1666464484
transform 1 0 116032 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1028
timestamp 1666464484
transform 1 0 116480 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_1031
timestamp 1666464484
transform 1 0 116816 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1095
timestamp 1666464484
transform 1 0 123984 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1099
timestamp 1666464484
transform 1 0 124432 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_1102
timestamp 1666464484
transform 1 0 124768 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1166
timestamp 1666464484
transform 1 0 131936 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1170
timestamp 1666464484
transform 1 0 132384 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_1173
timestamp 1666464484
transform 1 0 132720 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1237
timestamp 1666464484
transform 1 0 139888 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1241
timestamp 1666464484
transform 1 0 140336 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_1244
timestamp 1666464484
transform 1 0 140672 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1308
timestamp 1666464484
transform 1 0 147840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1312
timestamp 1666464484
transform 1 0 148288 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_1315
timestamp 1666464484
transform 1 0 148624 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1379
timestamp 1666464484
transform 1 0 155792 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1383
timestamp 1666464484
transform 1 0 156240 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_1386
timestamp 1666464484
transform 1 0 156576 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1450
timestamp 1666464484
transform 1 0 163744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1454
timestamp 1666464484
transform 1 0 164192 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_1457
timestamp 1666464484
transform 1 0 164528 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1521
timestamp 1666464484
transform 1 0 171696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1525
timestamp 1666464484
transform 1 0 172144 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_1528
timestamp 1666464484
transform 1 0 172480 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_1560
timestamp 1666464484
transform 1 0 176064 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1576
timestamp 1666464484
transform 1 0 177856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1580
timestamp 1666464484
transform 1 0 178304 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1666464484
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1666464484
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1666464484
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1666464484
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1666464484
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1666464484
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1666464484
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1666464484
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1666464484
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1666464484
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1666464484
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1666464484
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1666464484
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1666464484
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1666464484
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_357
timestamp 1666464484
transform 1 0 41328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_421
timestamp 1666464484
transform 1 0 48496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1666464484
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1666464484
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_492
timestamp 1666464484
transform 1 0 56448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1666464484
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_499
timestamp 1666464484
transform 1 0 57232 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_563
timestamp 1666464484
transform 1 0 64400 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_567
timestamp 1666464484
transform 1 0 64848 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_570
timestamp 1666464484
transform 1 0 65184 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_634
timestamp 1666464484
transform 1 0 72352 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_638
timestamp 1666464484
transform 1 0 72800 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_641
timestamp 1666464484
transform 1 0 73136 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_705
timestamp 1666464484
transform 1 0 80304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_709
timestamp 1666464484
transform 1 0 80752 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_712
timestamp 1666464484
transform 1 0 81088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_776
timestamp 1666464484
transform 1 0 88256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_780
timestamp 1666464484
transform 1 0 88704 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_783
timestamp 1666464484
transform 1 0 89040 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_847
timestamp 1666464484
transform 1 0 96208 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_851
timestamp 1666464484
transform 1 0 96656 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_854
timestamp 1666464484
transform 1 0 96992 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_918
timestamp 1666464484
transform 1 0 104160 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_922
timestamp 1666464484
transform 1 0 104608 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_925
timestamp 1666464484
transform 1 0 104944 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_989
timestamp 1666464484
transform 1 0 112112 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_993
timestamp 1666464484
transform 1 0 112560 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_996
timestamp 1666464484
transform 1 0 112896 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1060
timestamp 1666464484
transform 1 0 120064 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1064
timestamp 1666464484
transform 1 0 120512 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_1067
timestamp 1666464484
transform 1 0 120848 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1131
timestamp 1666464484
transform 1 0 128016 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1135
timestamp 1666464484
transform 1 0 128464 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_1138
timestamp 1666464484
transform 1 0 128800 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1202
timestamp 1666464484
transform 1 0 135968 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1206
timestamp 1666464484
transform 1 0 136416 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_1209
timestamp 1666464484
transform 1 0 136752 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1273
timestamp 1666464484
transform 1 0 143920 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1277
timestamp 1666464484
transform 1 0 144368 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_1280
timestamp 1666464484
transform 1 0 144704 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1344
timestamp 1666464484
transform 1 0 151872 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1348
timestamp 1666464484
transform 1 0 152320 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_1351
timestamp 1666464484
transform 1 0 152656 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1415
timestamp 1666464484
transform 1 0 159824 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1419
timestamp 1666464484
transform 1 0 160272 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_1422
timestamp 1666464484
transform 1 0 160608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1486
timestamp 1666464484
transform 1 0 167776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1490
timestamp 1666464484
transform 1 0 168224 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_1493
timestamp 1666464484
transform 1 0 168560 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_1557
timestamp 1666464484
transform 1 0 175728 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1561
timestamp 1666464484
transform 1 0 176176 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_1564
timestamp 1666464484
transform 1 0 176512 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1580
timestamp 1666464484
transform 1 0 178304 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_2
timestamp 1666464484
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1666464484
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1666464484
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1666464484
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1666464484
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1666464484
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1666464484
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1666464484
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1666464484
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1666464484
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1666464484
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1666464484
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1666464484
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1666464484
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1666464484
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1666464484
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1666464484
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_392
timestamp 1666464484
transform 1 0 45248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_456
timestamp 1666464484
transform 1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1666464484
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_463
timestamp 1666464484
transform 1 0 53200 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_527
timestamp 1666464484
transform 1 0 60368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 60816 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_534
timestamp 1666464484
transform 1 0 61152 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_598
timestamp 1666464484
transform 1 0 68320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_602
timestamp 1666464484
transform 1 0 68768 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_605
timestamp 1666464484
transform 1 0 69104 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_669
timestamp 1666464484
transform 1 0 76272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_673
timestamp 1666464484
transform 1 0 76720 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_676
timestamp 1666464484
transform 1 0 77056 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_740
timestamp 1666464484
transform 1 0 84224 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_744
timestamp 1666464484
transform 1 0 84672 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_747
timestamp 1666464484
transform 1 0 85008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_811
timestamp 1666464484
transform 1 0 92176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_815
timestamp 1666464484
transform 1 0 92624 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_818
timestamp 1666464484
transform 1 0 92960 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_882
timestamp 1666464484
transform 1 0 100128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_886
timestamp 1666464484
transform 1 0 100576 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_889
timestamp 1666464484
transform 1 0 100912 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_953
timestamp 1666464484
transform 1 0 108080 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_957
timestamp 1666464484
transform 1 0 108528 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_960
timestamp 1666464484
transform 1 0 108864 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1024
timestamp 1666464484
transform 1 0 116032 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1028
timestamp 1666464484
transform 1 0 116480 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_1031
timestamp 1666464484
transform 1 0 116816 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1095
timestamp 1666464484
transform 1 0 123984 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1099
timestamp 1666464484
transform 1 0 124432 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_1102
timestamp 1666464484
transform 1 0 124768 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1166
timestamp 1666464484
transform 1 0 131936 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1170
timestamp 1666464484
transform 1 0 132384 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_1173
timestamp 1666464484
transform 1 0 132720 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1237
timestamp 1666464484
transform 1 0 139888 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1241
timestamp 1666464484
transform 1 0 140336 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_1244
timestamp 1666464484
transform 1 0 140672 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1308
timestamp 1666464484
transform 1 0 147840 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1312
timestamp 1666464484
transform 1 0 148288 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_1315
timestamp 1666464484
transform 1 0 148624 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1379
timestamp 1666464484
transform 1 0 155792 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1383
timestamp 1666464484
transform 1 0 156240 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_1386
timestamp 1666464484
transform 1 0 156576 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1450
timestamp 1666464484
transform 1 0 163744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1454
timestamp 1666464484
transform 1 0 164192 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_1457
timestamp 1666464484
transform 1 0 164528 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1521
timestamp 1666464484
transform 1 0 171696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1525
timestamp 1666464484
transform 1 0 172144 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_1528
timestamp 1666464484
transform 1 0 172480 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_1560
timestamp 1666464484
transform 1 0 176064 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1576
timestamp 1666464484
transform 1 0 177856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1580
timestamp 1666464484
transform 1 0 178304 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1666464484
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1666464484
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1666464484
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1666464484
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1666464484
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1666464484
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1666464484
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1666464484
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1666464484
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1666464484
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1666464484
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1666464484
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1666464484
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1666464484
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1666464484
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_357
timestamp 1666464484
transform 1 0 41328 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_421
timestamp 1666464484
transform 1 0 48496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1666464484
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_428
timestamp 1666464484
transform 1 0 49280 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_492
timestamp 1666464484
transform 1 0 56448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1666464484
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_499
timestamp 1666464484
transform 1 0 57232 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_563
timestamp 1666464484
transform 1 0 64400 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_567
timestamp 1666464484
transform 1 0 64848 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_570
timestamp 1666464484
transform 1 0 65184 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_634
timestamp 1666464484
transform 1 0 72352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_638
timestamp 1666464484
transform 1 0 72800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_641
timestamp 1666464484
transform 1 0 73136 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_705
timestamp 1666464484
transform 1 0 80304 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_709
timestamp 1666464484
transform 1 0 80752 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_712
timestamp 1666464484
transform 1 0 81088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_776
timestamp 1666464484
transform 1 0 88256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_780
timestamp 1666464484
transform 1 0 88704 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_783
timestamp 1666464484
transform 1 0 89040 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_847
timestamp 1666464484
transform 1 0 96208 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_851
timestamp 1666464484
transform 1 0 96656 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_854
timestamp 1666464484
transform 1 0 96992 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_918
timestamp 1666464484
transform 1 0 104160 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_922
timestamp 1666464484
transform 1 0 104608 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_925
timestamp 1666464484
transform 1 0 104944 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_989
timestamp 1666464484
transform 1 0 112112 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_993
timestamp 1666464484
transform 1 0 112560 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_996
timestamp 1666464484
transform 1 0 112896 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1060
timestamp 1666464484
transform 1 0 120064 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1064
timestamp 1666464484
transform 1 0 120512 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_1067
timestamp 1666464484
transform 1 0 120848 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1131
timestamp 1666464484
transform 1 0 128016 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1135
timestamp 1666464484
transform 1 0 128464 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_1138
timestamp 1666464484
transform 1 0 128800 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1202
timestamp 1666464484
transform 1 0 135968 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1206
timestamp 1666464484
transform 1 0 136416 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_1209
timestamp 1666464484
transform 1 0 136752 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1273
timestamp 1666464484
transform 1 0 143920 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1277
timestamp 1666464484
transform 1 0 144368 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_1280
timestamp 1666464484
transform 1 0 144704 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1344
timestamp 1666464484
transform 1 0 151872 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1348
timestamp 1666464484
transform 1 0 152320 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_1351
timestamp 1666464484
transform 1 0 152656 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1415
timestamp 1666464484
transform 1 0 159824 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1419
timestamp 1666464484
transform 1 0 160272 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_1422
timestamp 1666464484
transform 1 0 160608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1486
timestamp 1666464484
transform 1 0 167776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1490
timestamp 1666464484
transform 1 0 168224 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_1493
timestamp 1666464484
transform 1 0 168560 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_1557
timestamp 1666464484
transform 1 0 175728 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1561
timestamp 1666464484
transform 1 0 176176 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_1564
timestamp 1666464484
transform 1 0 176512 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1580
timestamp 1666464484
transform 1 0 178304 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1666464484
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1666464484
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1666464484
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1666464484
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1666464484
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1666464484
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1666464484
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1666464484
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1666464484
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1666464484
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1666464484
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1666464484
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1666464484
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1666464484
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1666464484
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1666464484
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1666464484
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_392
timestamp 1666464484
transform 1 0 45248 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_456
timestamp 1666464484
transform 1 0 52416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1666464484
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_463
timestamp 1666464484
transform 1 0 53200 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_527
timestamp 1666464484
transform 1 0 60368 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 60816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_534
timestamp 1666464484
transform 1 0 61152 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_598
timestamp 1666464484
transform 1 0 68320 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_602
timestamp 1666464484
transform 1 0 68768 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_605
timestamp 1666464484
transform 1 0 69104 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_669
timestamp 1666464484
transform 1 0 76272 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_673
timestamp 1666464484
transform 1 0 76720 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_676
timestamp 1666464484
transform 1 0 77056 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_740
timestamp 1666464484
transform 1 0 84224 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_744
timestamp 1666464484
transform 1 0 84672 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_747
timestamp 1666464484
transform 1 0 85008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_811
timestamp 1666464484
transform 1 0 92176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_815
timestamp 1666464484
transform 1 0 92624 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_818
timestamp 1666464484
transform 1 0 92960 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_882
timestamp 1666464484
transform 1 0 100128 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_886
timestamp 1666464484
transform 1 0 100576 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_889
timestamp 1666464484
transform 1 0 100912 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_953
timestamp 1666464484
transform 1 0 108080 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_957
timestamp 1666464484
transform 1 0 108528 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_960
timestamp 1666464484
transform 1 0 108864 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1024
timestamp 1666464484
transform 1 0 116032 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1028
timestamp 1666464484
transform 1 0 116480 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_1031
timestamp 1666464484
transform 1 0 116816 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1095
timestamp 1666464484
transform 1 0 123984 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1099
timestamp 1666464484
transform 1 0 124432 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_1102
timestamp 1666464484
transform 1 0 124768 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1166
timestamp 1666464484
transform 1 0 131936 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1170
timestamp 1666464484
transform 1 0 132384 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_1173
timestamp 1666464484
transform 1 0 132720 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1237
timestamp 1666464484
transform 1 0 139888 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1241
timestamp 1666464484
transform 1 0 140336 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_1244
timestamp 1666464484
transform 1 0 140672 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1308
timestamp 1666464484
transform 1 0 147840 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1312
timestamp 1666464484
transform 1 0 148288 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_1315
timestamp 1666464484
transform 1 0 148624 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1379
timestamp 1666464484
transform 1 0 155792 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1383
timestamp 1666464484
transform 1 0 156240 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_1386
timestamp 1666464484
transform 1 0 156576 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1450
timestamp 1666464484
transform 1 0 163744 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1454
timestamp 1666464484
transform 1 0 164192 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_1457
timestamp 1666464484
transform 1 0 164528 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1521
timestamp 1666464484
transform 1 0 171696 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1525
timestamp 1666464484
transform 1 0 172144 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_1528
timestamp 1666464484
transform 1 0 172480 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_1560
timestamp 1666464484
transform 1 0 176064 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1576
timestamp 1666464484
transform 1 0 177856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1580
timestamp 1666464484
transform 1 0 178304 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1666464484
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1666464484
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1666464484
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1666464484
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1666464484
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1666464484
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1666464484
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1666464484
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1666464484
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1666464484
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1666464484
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1666464484
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1666464484
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1666464484
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1666464484
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_357
timestamp 1666464484
transform 1 0 41328 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_421
timestamp 1666464484
transform 1 0 48496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1666464484
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_428
timestamp 1666464484
transform 1 0 49280 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_492
timestamp 1666464484
transform 1 0 56448 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1666464484
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_499
timestamp 1666464484
transform 1 0 57232 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_563
timestamp 1666464484
transform 1 0 64400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_567
timestamp 1666464484
transform 1 0 64848 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_570
timestamp 1666464484
transform 1 0 65184 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_634
timestamp 1666464484
transform 1 0 72352 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_638
timestamp 1666464484
transform 1 0 72800 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_641
timestamp 1666464484
transform 1 0 73136 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_705
timestamp 1666464484
transform 1 0 80304 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_709
timestamp 1666464484
transform 1 0 80752 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_712
timestamp 1666464484
transform 1 0 81088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_776
timestamp 1666464484
transform 1 0 88256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_780
timestamp 1666464484
transform 1 0 88704 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_783
timestamp 1666464484
transform 1 0 89040 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_847
timestamp 1666464484
transform 1 0 96208 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_851
timestamp 1666464484
transform 1 0 96656 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_854
timestamp 1666464484
transform 1 0 96992 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_918
timestamp 1666464484
transform 1 0 104160 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_922
timestamp 1666464484
transform 1 0 104608 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_925
timestamp 1666464484
transform 1 0 104944 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_989
timestamp 1666464484
transform 1 0 112112 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_993
timestamp 1666464484
transform 1 0 112560 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_996
timestamp 1666464484
transform 1 0 112896 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1060
timestamp 1666464484
transform 1 0 120064 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1064
timestamp 1666464484
transform 1 0 120512 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_1067
timestamp 1666464484
transform 1 0 120848 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1131
timestamp 1666464484
transform 1 0 128016 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1135
timestamp 1666464484
transform 1 0 128464 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_1138
timestamp 1666464484
transform 1 0 128800 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1202
timestamp 1666464484
transform 1 0 135968 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1206
timestamp 1666464484
transform 1 0 136416 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_1209
timestamp 1666464484
transform 1 0 136752 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1273
timestamp 1666464484
transform 1 0 143920 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1277
timestamp 1666464484
transform 1 0 144368 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_1280
timestamp 1666464484
transform 1 0 144704 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1344
timestamp 1666464484
transform 1 0 151872 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1348
timestamp 1666464484
transform 1 0 152320 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_1351
timestamp 1666464484
transform 1 0 152656 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1415
timestamp 1666464484
transform 1 0 159824 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1419
timestamp 1666464484
transform 1 0 160272 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_1422
timestamp 1666464484
transform 1 0 160608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1486
timestamp 1666464484
transform 1 0 167776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1490
timestamp 1666464484
transform 1 0 168224 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_1493
timestamp 1666464484
transform 1 0 168560 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_1557
timestamp 1666464484
transform 1 0 175728 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1561
timestamp 1666464484
transform 1 0 176176 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_1564
timestamp 1666464484
transform 1 0 176512 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1580
timestamp 1666464484
transform 1 0 178304 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1666464484
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1666464484
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1666464484
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1666464484
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1666464484
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1666464484
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1666464484
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1666464484
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1666464484
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1666464484
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1666464484
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1666464484
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1666464484
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1666464484
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1666464484
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1666464484
transform 1 0 44464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1666464484
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_392
timestamp 1666464484
transform 1 0 45248 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_456
timestamp 1666464484
transform 1 0 52416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1666464484
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_463
timestamp 1666464484
transform 1 0 53200 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_527
timestamp 1666464484
transform 1 0 60368 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 60816 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_534
timestamp 1666464484
transform 1 0 61152 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_598
timestamp 1666464484
transform 1 0 68320 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_602
timestamp 1666464484
transform 1 0 68768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_605
timestamp 1666464484
transform 1 0 69104 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_669
timestamp 1666464484
transform 1 0 76272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_673
timestamp 1666464484
transform 1 0 76720 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_676
timestamp 1666464484
transform 1 0 77056 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_740
timestamp 1666464484
transform 1 0 84224 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_744
timestamp 1666464484
transform 1 0 84672 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_747
timestamp 1666464484
transform 1 0 85008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_811
timestamp 1666464484
transform 1 0 92176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_815
timestamp 1666464484
transform 1 0 92624 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_818
timestamp 1666464484
transform 1 0 92960 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_882
timestamp 1666464484
transform 1 0 100128 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_886
timestamp 1666464484
transform 1 0 100576 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_889
timestamp 1666464484
transform 1 0 100912 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_953
timestamp 1666464484
transform 1 0 108080 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_957
timestamp 1666464484
transform 1 0 108528 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_960
timestamp 1666464484
transform 1 0 108864 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1024
timestamp 1666464484
transform 1 0 116032 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1028
timestamp 1666464484
transform 1 0 116480 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_1031
timestamp 1666464484
transform 1 0 116816 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1095
timestamp 1666464484
transform 1 0 123984 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1099
timestamp 1666464484
transform 1 0 124432 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_1102
timestamp 1666464484
transform 1 0 124768 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1166
timestamp 1666464484
transform 1 0 131936 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1170
timestamp 1666464484
transform 1 0 132384 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_1173
timestamp 1666464484
transform 1 0 132720 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1237
timestamp 1666464484
transform 1 0 139888 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1241
timestamp 1666464484
transform 1 0 140336 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_1244
timestamp 1666464484
transform 1 0 140672 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1308
timestamp 1666464484
transform 1 0 147840 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1312
timestamp 1666464484
transform 1 0 148288 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_1315
timestamp 1666464484
transform 1 0 148624 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1379
timestamp 1666464484
transform 1 0 155792 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1383
timestamp 1666464484
transform 1 0 156240 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_1386
timestamp 1666464484
transform 1 0 156576 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1450
timestamp 1666464484
transform 1 0 163744 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1454
timestamp 1666464484
transform 1 0 164192 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_1457
timestamp 1666464484
transform 1 0 164528 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1521
timestamp 1666464484
transform 1 0 171696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1525
timestamp 1666464484
transform 1 0 172144 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_1528
timestamp 1666464484
transform 1 0 172480 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_1560
timestamp 1666464484
transform 1 0 176064 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1576
timestamp 1666464484
transform 1 0 177856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1580
timestamp 1666464484
transform 1 0 178304 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1666464484
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1666464484
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1666464484
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1666464484
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1666464484
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1666464484
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1666464484
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1666464484
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1666464484
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1666464484
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1666464484
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1666464484
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1666464484
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1666464484
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1666464484
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_357
timestamp 1666464484
transform 1 0 41328 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_421
timestamp 1666464484
transform 1 0 48496 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1666464484
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_428
timestamp 1666464484
transform 1 0 49280 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_492
timestamp 1666464484
transform 1 0 56448 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1666464484
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_499
timestamp 1666464484
transform 1 0 57232 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_563
timestamp 1666464484
transform 1 0 64400 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_567
timestamp 1666464484
transform 1 0 64848 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_570
timestamp 1666464484
transform 1 0 65184 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_634
timestamp 1666464484
transform 1 0 72352 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_638
timestamp 1666464484
transform 1 0 72800 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_641
timestamp 1666464484
transform 1 0 73136 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_705
timestamp 1666464484
transform 1 0 80304 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_709
timestamp 1666464484
transform 1 0 80752 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_712
timestamp 1666464484
transform 1 0 81088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_776
timestamp 1666464484
transform 1 0 88256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_780
timestamp 1666464484
transform 1 0 88704 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_783
timestamp 1666464484
transform 1 0 89040 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_847
timestamp 1666464484
transform 1 0 96208 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_851
timestamp 1666464484
transform 1 0 96656 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_854
timestamp 1666464484
transform 1 0 96992 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_918
timestamp 1666464484
transform 1 0 104160 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_922
timestamp 1666464484
transform 1 0 104608 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_925
timestamp 1666464484
transform 1 0 104944 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_989
timestamp 1666464484
transform 1 0 112112 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_993
timestamp 1666464484
transform 1 0 112560 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_996
timestamp 1666464484
transform 1 0 112896 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1060
timestamp 1666464484
transform 1 0 120064 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1064
timestamp 1666464484
transform 1 0 120512 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_1067
timestamp 1666464484
transform 1 0 120848 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1131
timestamp 1666464484
transform 1 0 128016 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1135
timestamp 1666464484
transform 1 0 128464 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_1138
timestamp 1666464484
transform 1 0 128800 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1202
timestamp 1666464484
transform 1 0 135968 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1206
timestamp 1666464484
transform 1 0 136416 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_1209
timestamp 1666464484
transform 1 0 136752 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1273
timestamp 1666464484
transform 1 0 143920 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1277
timestamp 1666464484
transform 1 0 144368 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_1280
timestamp 1666464484
transform 1 0 144704 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1344
timestamp 1666464484
transform 1 0 151872 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1348
timestamp 1666464484
transform 1 0 152320 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_1351
timestamp 1666464484
transform 1 0 152656 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1415
timestamp 1666464484
transform 1 0 159824 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1419
timestamp 1666464484
transform 1 0 160272 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_1422
timestamp 1666464484
transform 1 0 160608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1486
timestamp 1666464484
transform 1 0 167776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1490
timestamp 1666464484
transform 1 0 168224 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_1493
timestamp 1666464484
transform 1 0 168560 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_1557
timestamp 1666464484
transform 1 0 175728 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1561
timestamp 1666464484
transform 1 0 176176 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_1564
timestamp 1666464484
transform 1 0 176512 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1580
timestamp 1666464484
transform 1 0 178304 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1666464484
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1666464484
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1666464484
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1666464484
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1666464484
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1666464484
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1666464484
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1666464484
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1666464484
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1666464484
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1666464484
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1666464484
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1666464484
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1666464484
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1666464484
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_385
timestamp 1666464484
transform 1 0 44464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1666464484
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_392
timestamp 1666464484
transform 1 0 45248 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_456
timestamp 1666464484
transform 1 0 52416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1666464484
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_463
timestamp 1666464484
transform 1 0 53200 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_527
timestamp 1666464484
transform 1 0 60368 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_531
timestamp 1666464484
transform 1 0 60816 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_534
timestamp 1666464484
transform 1 0 61152 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_598
timestamp 1666464484
transform 1 0 68320 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_602
timestamp 1666464484
transform 1 0 68768 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_605
timestamp 1666464484
transform 1 0 69104 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_669
timestamp 1666464484
transform 1 0 76272 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_673
timestamp 1666464484
transform 1 0 76720 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_676
timestamp 1666464484
transform 1 0 77056 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_740
timestamp 1666464484
transform 1 0 84224 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_744
timestamp 1666464484
transform 1 0 84672 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_747
timestamp 1666464484
transform 1 0 85008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_811
timestamp 1666464484
transform 1 0 92176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_815
timestamp 1666464484
transform 1 0 92624 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_818
timestamp 1666464484
transform 1 0 92960 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_882
timestamp 1666464484
transform 1 0 100128 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_886
timestamp 1666464484
transform 1 0 100576 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_889
timestamp 1666464484
transform 1 0 100912 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_953
timestamp 1666464484
transform 1 0 108080 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_957
timestamp 1666464484
transform 1 0 108528 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_960
timestamp 1666464484
transform 1 0 108864 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1024
timestamp 1666464484
transform 1 0 116032 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1028
timestamp 1666464484
transform 1 0 116480 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_1031
timestamp 1666464484
transform 1 0 116816 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1095
timestamp 1666464484
transform 1 0 123984 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1099
timestamp 1666464484
transform 1 0 124432 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_1102
timestamp 1666464484
transform 1 0 124768 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1166
timestamp 1666464484
transform 1 0 131936 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1170
timestamp 1666464484
transform 1 0 132384 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_1173
timestamp 1666464484
transform 1 0 132720 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1237
timestamp 1666464484
transform 1 0 139888 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1241
timestamp 1666464484
transform 1 0 140336 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_1244
timestamp 1666464484
transform 1 0 140672 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1308
timestamp 1666464484
transform 1 0 147840 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1312
timestamp 1666464484
transform 1 0 148288 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_1315
timestamp 1666464484
transform 1 0 148624 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1379
timestamp 1666464484
transform 1 0 155792 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1383
timestamp 1666464484
transform 1 0 156240 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_1386
timestamp 1666464484
transform 1 0 156576 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1450
timestamp 1666464484
transform 1 0 163744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1454
timestamp 1666464484
transform 1 0 164192 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_1457
timestamp 1666464484
transform 1 0 164528 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1521
timestamp 1666464484
transform 1 0 171696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1525
timestamp 1666464484
transform 1 0 172144 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_1528
timestamp 1666464484
transform 1 0 172480 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_1560
timestamp 1666464484
transform 1 0 176064 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1576
timestamp 1666464484
transform 1 0 177856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1580
timestamp 1666464484
transform 1 0 178304 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1666464484
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1666464484
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1666464484
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1666464484
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1666464484
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1666464484
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1666464484
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1666464484
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1666464484
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1666464484
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1666464484
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1666464484
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1666464484
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1666464484
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1666464484
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_357
timestamp 1666464484
transform 1 0 41328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_421
timestamp 1666464484
transform 1 0 48496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1666464484
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_428
timestamp 1666464484
transform 1 0 49280 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_492
timestamp 1666464484
transform 1 0 56448 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1666464484
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_499
timestamp 1666464484
transform 1 0 57232 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_563
timestamp 1666464484
transform 1 0 64400 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_567
timestamp 1666464484
transform 1 0 64848 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_570
timestamp 1666464484
transform 1 0 65184 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_634
timestamp 1666464484
transform 1 0 72352 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_638
timestamp 1666464484
transform 1 0 72800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_641
timestamp 1666464484
transform 1 0 73136 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_705
timestamp 1666464484
transform 1 0 80304 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_709
timestamp 1666464484
transform 1 0 80752 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_712
timestamp 1666464484
transform 1 0 81088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_776
timestamp 1666464484
transform 1 0 88256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_780
timestamp 1666464484
transform 1 0 88704 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_783
timestamp 1666464484
transform 1 0 89040 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_847
timestamp 1666464484
transform 1 0 96208 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_851
timestamp 1666464484
transform 1 0 96656 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_854
timestamp 1666464484
transform 1 0 96992 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_918
timestamp 1666464484
transform 1 0 104160 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_922
timestamp 1666464484
transform 1 0 104608 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_925
timestamp 1666464484
transform 1 0 104944 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_989
timestamp 1666464484
transform 1 0 112112 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_993
timestamp 1666464484
transform 1 0 112560 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_996
timestamp 1666464484
transform 1 0 112896 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_1060
timestamp 1666464484
transform 1 0 120064 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1064
timestamp 1666464484
transform 1 0 120512 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_1067
timestamp 1666464484
transform 1 0 120848 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_1131
timestamp 1666464484
transform 1 0 128016 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1135
timestamp 1666464484
transform 1 0 128464 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_1138
timestamp 1666464484
transform 1 0 128800 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_1202
timestamp 1666464484
transform 1 0 135968 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1206
timestamp 1666464484
transform 1 0 136416 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_1209
timestamp 1666464484
transform 1 0 136752 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_1273
timestamp 1666464484
transform 1 0 143920 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1277
timestamp 1666464484
transform 1 0 144368 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_1280
timestamp 1666464484
transform 1 0 144704 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_1344
timestamp 1666464484
transform 1 0 151872 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1348
timestamp 1666464484
transform 1 0 152320 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_1351
timestamp 1666464484
transform 1 0 152656 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_1415
timestamp 1666464484
transform 1 0 159824 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1419
timestamp 1666464484
transform 1 0 160272 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_1422
timestamp 1666464484
transform 1 0 160608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_1486
timestamp 1666464484
transform 1 0 167776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1490
timestamp 1666464484
transform 1 0 168224 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_1493
timestamp 1666464484
transform 1 0 168560 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_1557
timestamp 1666464484
transform 1 0 175728 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1561
timestamp 1666464484
transform 1 0 176176 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_1564
timestamp 1666464484
transform 1 0 176512 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1580
timestamp 1666464484
transform 1 0 178304 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1666464484
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1666464484
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1666464484
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1666464484
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1666464484
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1666464484
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1666464484
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1666464484
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1666464484
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1666464484
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1666464484
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1666464484
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1666464484
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1666464484
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1666464484
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1666464484
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1666464484
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_392
timestamp 1666464484
transform 1 0 45248 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_456
timestamp 1666464484
transform 1 0 52416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1666464484
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_463
timestamp 1666464484
transform 1 0 53200 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_527
timestamp 1666464484
transform 1 0 60368 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 60816 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_534
timestamp 1666464484
transform 1 0 61152 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_598
timestamp 1666464484
transform 1 0 68320 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_602
timestamp 1666464484
transform 1 0 68768 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_605
timestamp 1666464484
transform 1 0 69104 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_669
timestamp 1666464484
transform 1 0 76272 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_673
timestamp 1666464484
transform 1 0 76720 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_676
timestamp 1666464484
transform 1 0 77056 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_740
timestamp 1666464484
transform 1 0 84224 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_744
timestamp 1666464484
transform 1 0 84672 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_747
timestamp 1666464484
transform 1 0 85008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_811
timestamp 1666464484
transform 1 0 92176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_815
timestamp 1666464484
transform 1 0 92624 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_818
timestamp 1666464484
transform 1 0 92960 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_882
timestamp 1666464484
transform 1 0 100128 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_886
timestamp 1666464484
transform 1 0 100576 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_889
timestamp 1666464484
transform 1 0 100912 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_953
timestamp 1666464484
transform 1 0 108080 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_957
timestamp 1666464484
transform 1 0 108528 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_960
timestamp 1666464484
transform 1 0 108864 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1024
timestamp 1666464484
transform 1 0 116032 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1028
timestamp 1666464484
transform 1 0 116480 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_1031
timestamp 1666464484
transform 1 0 116816 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1095
timestamp 1666464484
transform 1 0 123984 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1099
timestamp 1666464484
transform 1 0 124432 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_1102
timestamp 1666464484
transform 1 0 124768 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1166
timestamp 1666464484
transform 1 0 131936 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1170
timestamp 1666464484
transform 1 0 132384 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_1173
timestamp 1666464484
transform 1 0 132720 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1237
timestamp 1666464484
transform 1 0 139888 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1241
timestamp 1666464484
transform 1 0 140336 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_1244
timestamp 1666464484
transform 1 0 140672 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1308
timestamp 1666464484
transform 1 0 147840 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1312
timestamp 1666464484
transform 1 0 148288 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_1315
timestamp 1666464484
transform 1 0 148624 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1379
timestamp 1666464484
transform 1 0 155792 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1383
timestamp 1666464484
transform 1 0 156240 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_1386
timestamp 1666464484
transform 1 0 156576 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1450
timestamp 1666464484
transform 1 0 163744 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1454
timestamp 1666464484
transform 1 0 164192 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_1457
timestamp 1666464484
transform 1 0 164528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1521
timestamp 1666464484
transform 1 0 171696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1525
timestamp 1666464484
transform 1 0 172144 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_1528
timestamp 1666464484
transform 1 0 172480 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_1560
timestamp 1666464484
transform 1 0 176064 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1576
timestamp 1666464484
transform 1 0 177856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1580
timestamp 1666464484
transform 1 0 178304 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1666464484
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1666464484
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1666464484
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1666464484
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1666464484
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1666464484
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1666464484
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1666464484
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1666464484
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1666464484
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1666464484
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1666464484
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1666464484
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1666464484
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1666464484
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_357
timestamp 1666464484
transform 1 0 41328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_421
timestamp 1666464484
transform 1 0 48496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1666464484
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1666464484
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_492
timestamp 1666464484
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1666464484
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_499
timestamp 1666464484
transform 1 0 57232 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_563
timestamp 1666464484
transform 1 0 64400 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_567
timestamp 1666464484
transform 1 0 64848 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_570
timestamp 1666464484
transform 1 0 65184 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_634
timestamp 1666464484
transform 1 0 72352 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_638
timestamp 1666464484
transform 1 0 72800 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_641
timestamp 1666464484
transform 1 0 73136 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_705
timestamp 1666464484
transform 1 0 80304 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_709
timestamp 1666464484
transform 1 0 80752 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_712
timestamp 1666464484
transform 1 0 81088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_776
timestamp 1666464484
transform 1 0 88256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_780
timestamp 1666464484
transform 1 0 88704 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_783
timestamp 1666464484
transform 1 0 89040 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_847
timestamp 1666464484
transform 1 0 96208 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_851
timestamp 1666464484
transform 1 0 96656 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_854
timestamp 1666464484
transform 1 0 96992 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_918
timestamp 1666464484
transform 1 0 104160 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_922
timestamp 1666464484
transform 1 0 104608 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_925
timestamp 1666464484
transform 1 0 104944 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_989
timestamp 1666464484
transform 1 0 112112 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_993
timestamp 1666464484
transform 1 0 112560 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_996
timestamp 1666464484
transform 1 0 112896 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1060
timestamp 1666464484
transform 1 0 120064 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1064
timestamp 1666464484
transform 1 0 120512 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_1067
timestamp 1666464484
transform 1 0 120848 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1131
timestamp 1666464484
transform 1 0 128016 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1135
timestamp 1666464484
transform 1 0 128464 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_1138
timestamp 1666464484
transform 1 0 128800 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1202
timestamp 1666464484
transform 1 0 135968 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1206
timestamp 1666464484
transform 1 0 136416 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_1209
timestamp 1666464484
transform 1 0 136752 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1273
timestamp 1666464484
transform 1 0 143920 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1277
timestamp 1666464484
transform 1 0 144368 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_1280
timestamp 1666464484
transform 1 0 144704 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1344
timestamp 1666464484
transform 1 0 151872 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1348
timestamp 1666464484
transform 1 0 152320 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_1351
timestamp 1666464484
transform 1 0 152656 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1415
timestamp 1666464484
transform 1 0 159824 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1419
timestamp 1666464484
transform 1 0 160272 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_1422
timestamp 1666464484
transform 1 0 160608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1486
timestamp 1666464484
transform 1 0 167776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1490
timestamp 1666464484
transform 1 0 168224 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_1493
timestamp 1666464484
transform 1 0 168560 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1557
timestamp 1666464484
transform 1 0 175728 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1561
timestamp 1666464484
transform 1 0 176176 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_1564
timestamp 1666464484
transform 1 0 176512 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1580
timestamp 1666464484
transform 1 0 178304 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1666464484
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1666464484
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1666464484
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1666464484
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1666464484
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1666464484
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1666464484
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1666464484
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1666464484
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1666464484
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1666464484
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1666464484
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1666464484
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1666464484
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1666464484
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1666464484
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1666464484
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_392
timestamp 1666464484
transform 1 0 45248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_456
timestamp 1666464484
transform 1 0 52416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1666464484
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_463
timestamp 1666464484
transform 1 0 53200 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_527
timestamp 1666464484
transform 1 0 60368 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_531
timestamp 1666464484
transform 1 0 60816 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_534
timestamp 1666464484
transform 1 0 61152 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_598
timestamp 1666464484
transform 1 0 68320 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_602
timestamp 1666464484
transform 1 0 68768 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_605
timestamp 1666464484
transform 1 0 69104 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_669
timestamp 1666464484
transform 1 0 76272 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_673
timestamp 1666464484
transform 1 0 76720 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_676
timestamp 1666464484
transform 1 0 77056 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_740
timestamp 1666464484
transform 1 0 84224 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_744
timestamp 1666464484
transform 1 0 84672 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_747
timestamp 1666464484
transform 1 0 85008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_811
timestamp 1666464484
transform 1 0 92176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_815
timestamp 1666464484
transform 1 0 92624 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_818
timestamp 1666464484
transform 1 0 92960 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_882
timestamp 1666464484
transform 1 0 100128 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_886
timestamp 1666464484
transform 1 0 100576 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_889
timestamp 1666464484
transform 1 0 100912 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_953
timestamp 1666464484
transform 1 0 108080 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_957
timestamp 1666464484
transform 1 0 108528 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_960
timestamp 1666464484
transform 1 0 108864 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1024
timestamp 1666464484
transform 1 0 116032 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1028
timestamp 1666464484
transform 1 0 116480 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_1031
timestamp 1666464484
transform 1 0 116816 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1095
timestamp 1666464484
transform 1 0 123984 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1099
timestamp 1666464484
transform 1 0 124432 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_1102
timestamp 1666464484
transform 1 0 124768 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1166
timestamp 1666464484
transform 1 0 131936 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1170
timestamp 1666464484
transform 1 0 132384 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_1173
timestamp 1666464484
transform 1 0 132720 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1237
timestamp 1666464484
transform 1 0 139888 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1241
timestamp 1666464484
transform 1 0 140336 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_1244
timestamp 1666464484
transform 1 0 140672 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1308
timestamp 1666464484
transform 1 0 147840 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1312
timestamp 1666464484
transform 1 0 148288 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_1315
timestamp 1666464484
transform 1 0 148624 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1379
timestamp 1666464484
transform 1 0 155792 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1383
timestamp 1666464484
transform 1 0 156240 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_1386
timestamp 1666464484
transform 1 0 156576 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1450
timestamp 1666464484
transform 1 0 163744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1454
timestamp 1666464484
transform 1 0 164192 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_1457
timestamp 1666464484
transform 1 0 164528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1521
timestamp 1666464484
transform 1 0 171696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1525
timestamp 1666464484
transform 1 0 172144 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_1528
timestamp 1666464484
transform 1 0 172480 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_1560
timestamp 1666464484
transform 1 0 176064 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1576
timestamp 1666464484
transform 1 0 177856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1580
timestamp 1666464484
transform 1 0 178304 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1666464484
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1666464484
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1666464484
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1666464484
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1666464484
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1666464484
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1666464484
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1666464484
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1666464484
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1666464484
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1666464484
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1666464484
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1666464484
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1666464484
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1666464484
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1666464484
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_421
timestamp 1666464484
transform 1 0 48496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1666464484
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1666464484
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_492
timestamp 1666464484
transform 1 0 56448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1666464484
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_499
timestamp 1666464484
transform 1 0 57232 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_563
timestamp 1666464484
transform 1 0 64400 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_567
timestamp 1666464484
transform 1 0 64848 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_570
timestamp 1666464484
transform 1 0 65184 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_634
timestamp 1666464484
transform 1 0 72352 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_638
timestamp 1666464484
transform 1 0 72800 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_641
timestamp 1666464484
transform 1 0 73136 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_705
timestamp 1666464484
transform 1 0 80304 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_709
timestamp 1666464484
transform 1 0 80752 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_712
timestamp 1666464484
transform 1 0 81088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_776
timestamp 1666464484
transform 1 0 88256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_780
timestamp 1666464484
transform 1 0 88704 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_783
timestamp 1666464484
transform 1 0 89040 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_847
timestamp 1666464484
transform 1 0 96208 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_851
timestamp 1666464484
transform 1 0 96656 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_854
timestamp 1666464484
transform 1 0 96992 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_918
timestamp 1666464484
transform 1 0 104160 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_922
timestamp 1666464484
transform 1 0 104608 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_925
timestamp 1666464484
transform 1 0 104944 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_989
timestamp 1666464484
transform 1 0 112112 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_993
timestamp 1666464484
transform 1 0 112560 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_996
timestamp 1666464484
transform 1 0 112896 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_1060
timestamp 1666464484
transform 1 0 120064 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1064
timestamp 1666464484
transform 1 0 120512 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_1067
timestamp 1666464484
transform 1 0 120848 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_1131
timestamp 1666464484
transform 1 0 128016 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1135
timestamp 1666464484
transform 1 0 128464 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_1138
timestamp 1666464484
transform 1 0 128800 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_1202
timestamp 1666464484
transform 1 0 135968 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1206
timestamp 1666464484
transform 1 0 136416 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_1209
timestamp 1666464484
transform 1 0 136752 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_1273
timestamp 1666464484
transform 1 0 143920 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1277
timestamp 1666464484
transform 1 0 144368 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_1280
timestamp 1666464484
transform 1 0 144704 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_1344
timestamp 1666464484
transform 1 0 151872 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1348
timestamp 1666464484
transform 1 0 152320 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_1351
timestamp 1666464484
transform 1 0 152656 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_1415
timestamp 1666464484
transform 1 0 159824 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1419
timestamp 1666464484
transform 1 0 160272 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_1422
timestamp 1666464484
transform 1 0 160608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_1486
timestamp 1666464484
transform 1 0 167776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1490
timestamp 1666464484
transform 1 0 168224 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_1493
timestamp 1666464484
transform 1 0 168560 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_1557
timestamp 1666464484
transform 1 0 175728 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1561
timestamp 1666464484
transform 1 0 176176 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_1564
timestamp 1666464484
transform 1 0 176512 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1580
timestamp 1666464484
transform 1 0 178304 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1666464484
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1666464484
transform 1 0 5152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1666464484
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1666464484
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1666464484
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1666464484
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1666464484
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1666464484
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1666464484
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1666464484
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1666464484
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1666464484
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1666464484
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1666464484
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1666464484
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1666464484
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1666464484
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_392
timestamp 1666464484
transform 1 0 45248 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_456
timestamp 1666464484
transform 1 0 52416 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1666464484
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_463
timestamp 1666464484
transform 1 0 53200 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_527
timestamp 1666464484
transform 1 0 60368 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 60816 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_534
timestamp 1666464484
transform 1 0 61152 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_598
timestamp 1666464484
transform 1 0 68320 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_602
timestamp 1666464484
transform 1 0 68768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_605
timestamp 1666464484
transform 1 0 69104 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_669
timestamp 1666464484
transform 1 0 76272 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_673
timestamp 1666464484
transform 1 0 76720 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_676
timestamp 1666464484
transform 1 0 77056 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_740
timestamp 1666464484
transform 1 0 84224 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_744
timestamp 1666464484
transform 1 0 84672 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_747
timestamp 1666464484
transform 1 0 85008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_811
timestamp 1666464484
transform 1 0 92176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_815
timestamp 1666464484
transform 1 0 92624 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_818
timestamp 1666464484
transform 1 0 92960 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_882
timestamp 1666464484
transform 1 0 100128 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_886
timestamp 1666464484
transform 1 0 100576 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_889
timestamp 1666464484
transform 1 0 100912 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_953
timestamp 1666464484
transform 1 0 108080 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_957
timestamp 1666464484
transform 1 0 108528 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_960
timestamp 1666464484
transform 1 0 108864 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1024
timestamp 1666464484
transform 1 0 116032 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1028
timestamp 1666464484
transform 1 0 116480 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_1031
timestamp 1666464484
transform 1 0 116816 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1095
timestamp 1666464484
transform 1 0 123984 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1099
timestamp 1666464484
transform 1 0 124432 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_1102
timestamp 1666464484
transform 1 0 124768 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1166
timestamp 1666464484
transform 1 0 131936 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1170
timestamp 1666464484
transform 1 0 132384 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_1173
timestamp 1666464484
transform 1 0 132720 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1237
timestamp 1666464484
transform 1 0 139888 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1241
timestamp 1666464484
transform 1 0 140336 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_1244
timestamp 1666464484
transform 1 0 140672 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1308
timestamp 1666464484
transform 1 0 147840 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1312
timestamp 1666464484
transform 1 0 148288 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_1315
timestamp 1666464484
transform 1 0 148624 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1379
timestamp 1666464484
transform 1 0 155792 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1383
timestamp 1666464484
transform 1 0 156240 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_1386
timestamp 1666464484
transform 1 0 156576 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1450
timestamp 1666464484
transform 1 0 163744 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1454
timestamp 1666464484
transform 1 0 164192 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_1457
timestamp 1666464484
transform 1 0 164528 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1521
timestamp 1666464484
transform 1 0 171696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1525
timestamp 1666464484
transform 1 0 172144 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_1528
timestamp 1666464484
transform 1 0 172480 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_1560
timestamp 1666464484
transform 1 0 176064 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1576
timestamp 1666464484
transform 1 0 177856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1580
timestamp 1666464484
transform 1 0 178304 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1666464484
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1666464484
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_70
timestamp 1666464484
transform 1 0 9184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_73
timestamp 1666464484
transform 1 0 9520 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_137
timestamp 1666464484
transform 1 0 16688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1666464484
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1666464484
transform 1 0 17472 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_208
timestamp 1666464484
transform 1 0 24640 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1666464484
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1666464484
transform 1 0 25424 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_279
timestamp 1666464484
transform 1 0 32592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1666464484
transform 1 0 33040 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1666464484
transform 1 0 33376 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1666464484
transform 1 0 40544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1666464484
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_357
timestamp 1666464484
transform 1 0 41328 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_421
timestamp 1666464484
transform 1 0 48496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_425
timestamp 1666464484
transform 1 0 48944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_428
timestamp 1666464484
transform 1 0 49280 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_492
timestamp 1666464484
transform 1 0 56448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1666464484
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_499
timestamp 1666464484
transform 1 0 57232 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_563
timestamp 1666464484
transform 1 0 64400 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_567
timestamp 1666464484
transform 1 0 64848 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_570
timestamp 1666464484
transform 1 0 65184 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_634
timestamp 1666464484
transform 1 0 72352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_638
timestamp 1666464484
transform 1 0 72800 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_641
timestamp 1666464484
transform 1 0 73136 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_705
timestamp 1666464484
transform 1 0 80304 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_709
timestamp 1666464484
transform 1 0 80752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_712
timestamp 1666464484
transform 1 0 81088 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_776
timestamp 1666464484
transform 1 0 88256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_780
timestamp 1666464484
transform 1 0 88704 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_783
timestamp 1666464484
transform 1 0 89040 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_847
timestamp 1666464484
transform 1 0 96208 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_851
timestamp 1666464484
transform 1 0 96656 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_854
timestamp 1666464484
transform 1 0 96992 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_918
timestamp 1666464484
transform 1 0 104160 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_922
timestamp 1666464484
transform 1 0 104608 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_925
timestamp 1666464484
transform 1 0 104944 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_989
timestamp 1666464484
transform 1 0 112112 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_993
timestamp 1666464484
transform 1 0 112560 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_996
timestamp 1666464484
transform 1 0 112896 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1060
timestamp 1666464484
transform 1 0 120064 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1064
timestamp 1666464484
transform 1 0 120512 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_1067
timestamp 1666464484
transform 1 0 120848 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1131
timestamp 1666464484
transform 1 0 128016 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1135
timestamp 1666464484
transform 1 0 128464 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_1138
timestamp 1666464484
transform 1 0 128800 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1202
timestamp 1666464484
transform 1 0 135968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1206
timestamp 1666464484
transform 1 0 136416 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_1209
timestamp 1666464484
transform 1 0 136752 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1273
timestamp 1666464484
transform 1 0 143920 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1277
timestamp 1666464484
transform 1 0 144368 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_1280
timestamp 1666464484
transform 1 0 144704 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1344
timestamp 1666464484
transform 1 0 151872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1348
timestamp 1666464484
transform 1 0 152320 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_1351
timestamp 1666464484
transform 1 0 152656 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1415
timestamp 1666464484
transform 1 0 159824 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1419
timestamp 1666464484
transform 1 0 160272 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_1422
timestamp 1666464484
transform 1 0 160608 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1486
timestamp 1666464484
transform 1 0 167776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1490
timestamp 1666464484
transform 1 0 168224 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_1493
timestamp 1666464484
transform 1 0 168560 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_1557
timestamp 1666464484
transform 1 0 175728 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1561
timestamp 1666464484
transform 1 0 176176 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_1564
timestamp 1666464484
transform 1 0 176512 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1580
timestamp 1666464484
transform 1 0 178304 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_2
timestamp 1666464484
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1666464484
transform 1 0 5152 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1666464484
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1666464484
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1666464484
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_108
timestamp 1666464484
transform 1 0 13440 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_172
timestamp 1666464484
transform 1 0 20608 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1666464484
transform 1 0 21056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1666464484
transform 1 0 21392 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_243
timestamp 1666464484
transform 1 0 28560 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1666464484
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1666464484
transform 1 0 29344 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_314
timestamp 1666464484
transform 1 0 36512 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1666464484
transform 1 0 36960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_321
timestamp 1666464484
transform 1 0 37296 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_385
timestamp 1666464484
transform 1 0 44464 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1666464484
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_392
timestamp 1666464484
transform 1 0 45248 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_456
timestamp 1666464484
transform 1 0 52416 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1666464484
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_463
timestamp 1666464484
transform 1 0 53200 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_527
timestamp 1666464484
transform 1 0 60368 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_531
timestamp 1666464484
transform 1 0 60816 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_534
timestamp 1666464484
transform 1 0 61152 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_598
timestamp 1666464484
transform 1 0 68320 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_602
timestamp 1666464484
transform 1 0 68768 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_605
timestamp 1666464484
transform 1 0 69104 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_669
timestamp 1666464484
transform 1 0 76272 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_673
timestamp 1666464484
transform 1 0 76720 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_676
timestamp 1666464484
transform 1 0 77056 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_740
timestamp 1666464484
transform 1 0 84224 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_744
timestamp 1666464484
transform 1 0 84672 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_747
timestamp 1666464484
transform 1 0 85008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_811
timestamp 1666464484
transform 1 0 92176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_815
timestamp 1666464484
transform 1 0 92624 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_818
timestamp 1666464484
transform 1 0 92960 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_882
timestamp 1666464484
transform 1 0 100128 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_886
timestamp 1666464484
transform 1 0 100576 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_889
timestamp 1666464484
transform 1 0 100912 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_953
timestamp 1666464484
transform 1 0 108080 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_957
timestamp 1666464484
transform 1 0 108528 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_960
timestamp 1666464484
transform 1 0 108864 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1024
timestamp 1666464484
transform 1 0 116032 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1028
timestamp 1666464484
transform 1 0 116480 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_1031
timestamp 1666464484
transform 1 0 116816 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1095
timestamp 1666464484
transform 1 0 123984 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1099
timestamp 1666464484
transform 1 0 124432 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_1102
timestamp 1666464484
transform 1 0 124768 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1166
timestamp 1666464484
transform 1 0 131936 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1170
timestamp 1666464484
transform 1 0 132384 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_1173
timestamp 1666464484
transform 1 0 132720 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1237
timestamp 1666464484
transform 1 0 139888 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1241
timestamp 1666464484
transform 1 0 140336 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_1244
timestamp 1666464484
transform 1 0 140672 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1308
timestamp 1666464484
transform 1 0 147840 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1312
timestamp 1666464484
transform 1 0 148288 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_1315
timestamp 1666464484
transform 1 0 148624 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1379
timestamp 1666464484
transform 1 0 155792 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1383
timestamp 1666464484
transform 1 0 156240 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_1386
timestamp 1666464484
transform 1 0 156576 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1450
timestamp 1666464484
transform 1 0 163744 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1454
timestamp 1666464484
transform 1 0 164192 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_1457
timestamp 1666464484
transform 1 0 164528 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1521
timestamp 1666464484
transform 1 0 171696 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1525
timestamp 1666464484
transform 1 0 172144 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_1528
timestamp 1666464484
transform 1 0 172480 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_1560
timestamp 1666464484
transform 1 0 176064 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1576
timestamp 1666464484
transform 1 0 177856 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1580
timestamp 1666464484
transform 1 0 178304 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_2
timestamp 1666464484
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_66
timestamp 1666464484
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_70
timestamp 1666464484
transform 1 0 9184 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_73
timestamp 1666464484
transform 1 0 9520 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_137
timestamp 1666464484
transform 1 0 16688 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_141
timestamp 1666464484
transform 1 0 17136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1666464484
transform 1 0 17472 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_208
timestamp 1666464484
transform 1 0 24640 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1666464484
transform 1 0 25088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1666464484
transform 1 0 25424 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_279
timestamp 1666464484
transform 1 0 32592 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1666464484
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1666464484
transform 1 0 33376 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_350
timestamp 1666464484
transform 1 0 40544 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1666464484
transform 1 0 40992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_357
timestamp 1666464484
transform 1 0 41328 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_421
timestamp 1666464484
transform 1 0 48496 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_425
timestamp 1666464484
transform 1 0 48944 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_428
timestamp 1666464484
transform 1 0 49280 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_492
timestamp 1666464484
transform 1 0 56448 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_496
timestamp 1666464484
transform 1 0 56896 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_499
timestamp 1666464484
transform 1 0 57232 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_563
timestamp 1666464484
transform 1 0 64400 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_567
timestamp 1666464484
transform 1 0 64848 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_570
timestamp 1666464484
transform 1 0 65184 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_634
timestamp 1666464484
transform 1 0 72352 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_638
timestamp 1666464484
transform 1 0 72800 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_641
timestamp 1666464484
transform 1 0 73136 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_705
timestamp 1666464484
transform 1 0 80304 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_709
timestamp 1666464484
transform 1 0 80752 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_712
timestamp 1666464484
transform 1 0 81088 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_776
timestamp 1666464484
transform 1 0 88256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_780
timestamp 1666464484
transform 1 0 88704 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_783
timestamp 1666464484
transform 1 0 89040 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_847
timestamp 1666464484
transform 1 0 96208 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_851
timestamp 1666464484
transform 1 0 96656 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_854
timestamp 1666464484
transform 1 0 96992 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_918
timestamp 1666464484
transform 1 0 104160 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_922
timestamp 1666464484
transform 1 0 104608 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_925
timestamp 1666464484
transform 1 0 104944 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_989
timestamp 1666464484
transform 1 0 112112 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_993
timestamp 1666464484
transform 1 0 112560 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_996
timestamp 1666464484
transform 1 0 112896 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1060
timestamp 1666464484
transform 1 0 120064 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1064
timestamp 1666464484
transform 1 0 120512 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_1067
timestamp 1666464484
transform 1 0 120848 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1131
timestamp 1666464484
transform 1 0 128016 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1135
timestamp 1666464484
transform 1 0 128464 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_1138
timestamp 1666464484
transform 1 0 128800 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1202
timestamp 1666464484
transform 1 0 135968 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1206
timestamp 1666464484
transform 1 0 136416 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_1209
timestamp 1666464484
transform 1 0 136752 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1273
timestamp 1666464484
transform 1 0 143920 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1277
timestamp 1666464484
transform 1 0 144368 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_1280
timestamp 1666464484
transform 1 0 144704 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1344
timestamp 1666464484
transform 1 0 151872 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1348
timestamp 1666464484
transform 1 0 152320 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_1351
timestamp 1666464484
transform 1 0 152656 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1415
timestamp 1666464484
transform 1 0 159824 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1419
timestamp 1666464484
transform 1 0 160272 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_1422
timestamp 1666464484
transform 1 0 160608 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1486
timestamp 1666464484
transform 1 0 167776 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1490
timestamp 1666464484
transform 1 0 168224 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_1493
timestamp 1666464484
transform 1 0 168560 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1557
timestamp 1666464484
transform 1 0 175728 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1561
timestamp 1666464484
transform 1 0 176176 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_1564
timestamp 1666464484
transform 1 0 176512 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1580
timestamp 1666464484
transform 1 0 178304 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_2
timestamp 1666464484
transform 1 0 1568 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_34
timestamp 1666464484
transform 1 0 5152 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_37
timestamp 1666464484
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_101
timestamp 1666464484
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1666464484
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_108
timestamp 1666464484
transform 1 0 13440 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_172
timestamp 1666464484
transform 1 0 20608 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1666464484
transform 1 0 21056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1666464484
transform 1 0 21392 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_243
timestamp 1666464484
transform 1 0 28560 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1666464484
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1666464484
transform 1 0 29344 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_314
timestamp 1666464484
transform 1 0 36512 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1666464484
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1666464484
transform 1 0 37296 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_385
timestamp 1666464484
transform 1 0 44464 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1666464484
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_392
timestamp 1666464484
transform 1 0 45248 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_456
timestamp 1666464484
transform 1 0 52416 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1666464484
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_463
timestamp 1666464484
transform 1 0 53200 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_527
timestamp 1666464484
transform 1 0 60368 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_531
timestamp 1666464484
transform 1 0 60816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_534
timestamp 1666464484
transform 1 0 61152 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_598
timestamp 1666464484
transform 1 0 68320 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_602
timestamp 1666464484
transform 1 0 68768 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_605
timestamp 1666464484
transform 1 0 69104 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_669
timestamp 1666464484
transform 1 0 76272 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_673
timestamp 1666464484
transform 1 0 76720 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_676
timestamp 1666464484
transform 1 0 77056 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_740
timestamp 1666464484
transform 1 0 84224 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_744
timestamp 1666464484
transform 1 0 84672 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_747
timestamp 1666464484
transform 1 0 85008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_811
timestamp 1666464484
transform 1 0 92176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_815
timestamp 1666464484
transform 1 0 92624 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_818
timestamp 1666464484
transform 1 0 92960 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_882
timestamp 1666464484
transform 1 0 100128 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_886
timestamp 1666464484
transform 1 0 100576 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_889
timestamp 1666464484
transform 1 0 100912 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_953
timestamp 1666464484
transform 1 0 108080 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_957
timestamp 1666464484
transform 1 0 108528 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_960
timestamp 1666464484
transform 1 0 108864 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1024
timestamp 1666464484
transform 1 0 116032 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1028
timestamp 1666464484
transform 1 0 116480 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_1031
timestamp 1666464484
transform 1 0 116816 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1095
timestamp 1666464484
transform 1 0 123984 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1099
timestamp 1666464484
transform 1 0 124432 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_1102
timestamp 1666464484
transform 1 0 124768 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1166
timestamp 1666464484
transform 1 0 131936 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1170
timestamp 1666464484
transform 1 0 132384 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_1173
timestamp 1666464484
transform 1 0 132720 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1237
timestamp 1666464484
transform 1 0 139888 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1241
timestamp 1666464484
transform 1 0 140336 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_1244
timestamp 1666464484
transform 1 0 140672 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1308
timestamp 1666464484
transform 1 0 147840 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1312
timestamp 1666464484
transform 1 0 148288 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_1315
timestamp 1666464484
transform 1 0 148624 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1379
timestamp 1666464484
transform 1 0 155792 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1383
timestamp 1666464484
transform 1 0 156240 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_1386
timestamp 1666464484
transform 1 0 156576 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1450
timestamp 1666464484
transform 1 0 163744 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1454
timestamp 1666464484
transform 1 0 164192 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_1457
timestamp 1666464484
transform 1 0 164528 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1521
timestamp 1666464484
transform 1 0 171696 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1525
timestamp 1666464484
transform 1 0 172144 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_1528
timestamp 1666464484
transform 1 0 172480 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_1560
timestamp 1666464484
transform 1 0 176064 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1576
timestamp 1666464484
transform 1 0 177856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1580
timestamp 1666464484
transform 1 0 178304 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_2
timestamp 1666464484
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_66
timestamp 1666464484
transform 1 0 8736 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_70
timestamp 1666464484
transform 1 0 9184 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_73
timestamp 1666464484
transform 1 0 9520 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_137
timestamp 1666464484
transform 1 0 16688 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1666464484
transform 1 0 17136 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_144
timestamp 1666464484
transform 1 0 17472 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_208
timestamp 1666464484
transform 1 0 24640 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1666464484
transform 1 0 25088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1666464484
transform 1 0 25424 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_279
timestamp 1666464484
transform 1 0 32592 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1666464484
transform 1 0 33040 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1666464484
transform 1 0 33376 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_350
timestamp 1666464484
transform 1 0 40544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1666464484
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_357
timestamp 1666464484
transform 1 0 41328 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_421
timestamp 1666464484
transform 1 0 48496 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_425
timestamp 1666464484
transform 1 0 48944 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_428
timestamp 1666464484
transform 1 0 49280 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_492
timestamp 1666464484
transform 1 0 56448 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_496
timestamp 1666464484
transform 1 0 56896 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_499
timestamp 1666464484
transform 1 0 57232 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_563
timestamp 1666464484
transform 1 0 64400 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_567
timestamp 1666464484
transform 1 0 64848 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_570
timestamp 1666464484
transform 1 0 65184 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_634
timestamp 1666464484
transform 1 0 72352 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_638
timestamp 1666464484
transform 1 0 72800 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_641
timestamp 1666464484
transform 1 0 73136 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_705
timestamp 1666464484
transform 1 0 80304 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_709
timestamp 1666464484
transform 1 0 80752 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_712
timestamp 1666464484
transform 1 0 81088 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_776
timestamp 1666464484
transform 1 0 88256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_780
timestamp 1666464484
transform 1 0 88704 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_783
timestamp 1666464484
transform 1 0 89040 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_847
timestamp 1666464484
transform 1 0 96208 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_851
timestamp 1666464484
transform 1 0 96656 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_854
timestamp 1666464484
transform 1 0 96992 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_918
timestamp 1666464484
transform 1 0 104160 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_922
timestamp 1666464484
transform 1 0 104608 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_925
timestamp 1666464484
transform 1 0 104944 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_989
timestamp 1666464484
transform 1 0 112112 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_993
timestamp 1666464484
transform 1 0 112560 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_996
timestamp 1666464484
transform 1 0 112896 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1060
timestamp 1666464484
transform 1 0 120064 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1064
timestamp 1666464484
transform 1 0 120512 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_1067
timestamp 1666464484
transform 1 0 120848 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1131
timestamp 1666464484
transform 1 0 128016 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1135
timestamp 1666464484
transform 1 0 128464 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_1138
timestamp 1666464484
transform 1 0 128800 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1202
timestamp 1666464484
transform 1 0 135968 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1206
timestamp 1666464484
transform 1 0 136416 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_1209
timestamp 1666464484
transform 1 0 136752 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1273
timestamp 1666464484
transform 1 0 143920 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1277
timestamp 1666464484
transform 1 0 144368 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_1280
timestamp 1666464484
transform 1 0 144704 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1344
timestamp 1666464484
transform 1 0 151872 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1348
timestamp 1666464484
transform 1 0 152320 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_1351
timestamp 1666464484
transform 1 0 152656 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1415
timestamp 1666464484
transform 1 0 159824 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1419
timestamp 1666464484
transform 1 0 160272 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_1422
timestamp 1666464484
transform 1 0 160608 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1486
timestamp 1666464484
transform 1 0 167776 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1490
timestamp 1666464484
transform 1 0 168224 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_1493
timestamp 1666464484
transform 1 0 168560 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1557
timestamp 1666464484
transform 1 0 175728 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1561
timestamp 1666464484
transform 1 0 176176 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_1564
timestamp 1666464484
transform 1 0 176512 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1580
timestamp 1666464484
transform 1 0 178304 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_2
timestamp 1666464484
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_34
timestamp 1666464484
transform 1 0 5152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_37
timestamp 1666464484
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_101
timestamp 1666464484
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1666464484
transform 1 0 13104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_108
timestamp 1666464484
transform 1 0 13440 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_172
timestamp 1666464484
transform 1 0 20608 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1666464484
transform 1 0 21056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_179
timestamp 1666464484
transform 1 0 21392 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_243
timestamp 1666464484
transform 1 0 28560 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1666464484
transform 1 0 29008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1666464484
transform 1 0 29344 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_314
timestamp 1666464484
transform 1 0 36512 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1666464484
transform 1 0 36960 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1666464484
transform 1 0 37296 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_385
timestamp 1666464484
transform 1 0 44464 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1666464484
transform 1 0 44912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_392
timestamp 1666464484
transform 1 0 45248 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_456
timestamp 1666464484
transform 1 0 52416 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_460
timestamp 1666464484
transform 1 0 52864 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_463
timestamp 1666464484
transform 1 0 53200 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_527
timestamp 1666464484
transform 1 0 60368 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 60816 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_534
timestamp 1666464484
transform 1 0 61152 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_598
timestamp 1666464484
transform 1 0 68320 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_602
timestamp 1666464484
transform 1 0 68768 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_605
timestamp 1666464484
transform 1 0 69104 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_669
timestamp 1666464484
transform 1 0 76272 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_673
timestamp 1666464484
transform 1 0 76720 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_676
timestamp 1666464484
transform 1 0 77056 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_740
timestamp 1666464484
transform 1 0 84224 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_744
timestamp 1666464484
transform 1 0 84672 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_747
timestamp 1666464484
transform 1 0 85008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_811
timestamp 1666464484
transform 1 0 92176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_815
timestamp 1666464484
transform 1 0 92624 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_818
timestamp 1666464484
transform 1 0 92960 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_882
timestamp 1666464484
transform 1 0 100128 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_886
timestamp 1666464484
transform 1 0 100576 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_889
timestamp 1666464484
transform 1 0 100912 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_953
timestamp 1666464484
transform 1 0 108080 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_957
timestamp 1666464484
transform 1 0 108528 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_960
timestamp 1666464484
transform 1 0 108864 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1024
timestamp 1666464484
transform 1 0 116032 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1028
timestamp 1666464484
transform 1 0 116480 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_1031
timestamp 1666464484
transform 1 0 116816 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1095
timestamp 1666464484
transform 1 0 123984 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1099
timestamp 1666464484
transform 1 0 124432 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_1102
timestamp 1666464484
transform 1 0 124768 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1166
timestamp 1666464484
transform 1 0 131936 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1170
timestamp 1666464484
transform 1 0 132384 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_1173
timestamp 1666464484
transform 1 0 132720 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1237
timestamp 1666464484
transform 1 0 139888 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1241
timestamp 1666464484
transform 1 0 140336 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_1244
timestamp 1666464484
transform 1 0 140672 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1308
timestamp 1666464484
transform 1 0 147840 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1312
timestamp 1666464484
transform 1 0 148288 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_1315
timestamp 1666464484
transform 1 0 148624 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1379
timestamp 1666464484
transform 1 0 155792 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1383
timestamp 1666464484
transform 1 0 156240 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_1386
timestamp 1666464484
transform 1 0 156576 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1450
timestamp 1666464484
transform 1 0 163744 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1454
timestamp 1666464484
transform 1 0 164192 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_1457
timestamp 1666464484
transform 1 0 164528 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1521
timestamp 1666464484
transform 1 0 171696 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1525
timestamp 1666464484
transform 1 0 172144 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_1528
timestamp 1666464484
transform 1 0 172480 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_1560
timestamp 1666464484
transform 1 0 176064 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1576
timestamp 1666464484
transform 1 0 177856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1580
timestamp 1666464484
transform 1 0 178304 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_2
timestamp 1666464484
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_66
timestamp 1666464484
transform 1 0 8736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_70
timestamp 1666464484
transform 1 0 9184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_73
timestamp 1666464484
transform 1 0 9520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_137
timestamp 1666464484
transform 1 0 16688 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1666464484
transform 1 0 17136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_144
timestamp 1666464484
transform 1 0 17472 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_208
timestamp 1666464484
transform 1 0 24640 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_212
timestamp 1666464484
transform 1 0 25088 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_215
timestamp 1666464484
transform 1 0 25424 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_279
timestamp 1666464484
transform 1 0 32592 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_283
timestamp 1666464484
transform 1 0 33040 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1666464484
transform 1 0 33376 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_350
timestamp 1666464484
transform 1 0 40544 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1666464484
transform 1 0 40992 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_357
timestamp 1666464484
transform 1 0 41328 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_421
timestamp 1666464484
transform 1 0 48496 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_425
timestamp 1666464484
transform 1 0 48944 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_428
timestamp 1666464484
transform 1 0 49280 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_492
timestamp 1666464484
transform 1 0 56448 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_496
timestamp 1666464484
transform 1 0 56896 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_499
timestamp 1666464484
transform 1 0 57232 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_563
timestamp 1666464484
transform 1 0 64400 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_567
timestamp 1666464484
transform 1 0 64848 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_570
timestamp 1666464484
transform 1 0 65184 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_634
timestamp 1666464484
transform 1 0 72352 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_638
timestamp 1666464484
transform 1 0 72800 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_641
timestamp 1666464484
transform 1 0 73136 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_705
timestamp 1666464484
transform 1 0 80304 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_709
timestamp 1666464484
transform 1 0 80752 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_712
timestamp 1666464484
transform 1 0 81088 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_776
timestamp 1666464484
transform 1 0 88256 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_780
timestamp 1666464484
transform 1 0 88704 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_783
timestamp 1666464484
transform 1 0 89040 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_847
timestamp 1666464484
transform 1 0 96208 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_851
timestamp 1666464484
transform 1 0 96656 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_854
timestamp 1666464484
transform 1 0 96992 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_918
timestamp 1666464484
transform 1 0 104160 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_922
timestamp 1666464484
transform 1 0 104608 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_925
timestamp 1666464484
transform 1 0 104944 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_989
timestamp 1666464484
transform 1 0 112112 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_993
timestamp 1666464484
transform 1 0 112560 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_996
timestamp 1666464484
transform 1 0 112896 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1060
timestamp 1666464484
transform 1 0 120064 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1064
timestamp 1666464484
transform 1 0 120512 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_1067
timestamp 1666464484
transform 1 0 120848 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1131
timestamp 1666464484
transform 1 0 128016 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1135
timestamp 1666464484
transform 1 0 128464 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_1138
timestamp 1666464484
transform 1 0 128800 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1202
timestamp 1666464484
transform 1 0 135968 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1206
timestamp 1666464484
transform 1 0 136416 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_1209
timestamp 1666464484
transform 1 0 136752 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1273
timestamp 1666464484
transform 1 0 143920 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1277
timestamp 1666464484
transform 1 0 144368 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_1280
timestamp 1666464484
transform 1 0 144704 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1344
timestamp 1666464484
transform 1 0 151872 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1348
timestamp 1666464484
transform 1 0 152320 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_1351
timestamp 1666464484
transform 1 0 152656 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1415
timestamp 1666464484
transform 1 0 159824 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1419
timestamp 1666464484
transform 1 0 160272 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_1422
timestamp 1666464484
transform 1 0 160608 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1486
timestamp 1666464484
transform 1 0 167776 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1490
timestamp 1666464484
transform 1 0 168224 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_1493
timestamp 1666464484
transform 1 0 168560 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1557
timestamp 1666464484
transform 1 0 175728 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1561
timestamp 1666464484
transform 1 0 176176 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_1564
timestamp 1666464484
transform 1 0 176512 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1580
timestamp 1666464484
transform 1 0 178304 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_2
timestamp 1666464484
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_34
timestamp 1666464484
transform 1 0 5152 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_37
timestamp 1666464484
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_101
timestamp 1666464484
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1666464484
transform 1 0 13104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_108
timestamp 1666464484
transform 1 0 13440 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_172
timestamp 1666464484
transform 1 0 20608 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_176
timestamp 1666464484
transform 1 0 21056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_179
timestamp 1666464484
transform 1 0 21392 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_243
timestamp 1666464484
transform 1 0 28560 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_247
timestamp 1666464484
transform 1 0 29008 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1666464484
transform 1 0 29344 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_314
timestamp 1666464484
transform 1 0 36512 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1666464484
transform 1 0 36960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1666464484
transform 1 0 37296 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_385
timestamp 1666464484
transform 1 0 44464 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1666464484
transform 1 0 44912 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_392
timestamp 1666464484
transform 1 0 45248 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_456
timestamp 1666464484
transform 1 0 52416 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_460
timestamp 1666464484
transform 1 0 52864 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_463
timestamp 1666464484
transform 1 0 53200 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_527
timestamp 1666464484
transform 1 0 60368 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_531
timestamp 1666464484
transform 1 0 60816 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_534
timestamp 1666464484
transform 1 0 61152 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_598
timestamp 1666464484
transform 1 0 68320 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_602
timestamp 1666464484
transform 1 0 68768 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_605
timestamp 1666464484
transform 1 0 69104 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_669
timestamp 1666464484
transform 1 0 76272 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_673
timestamp 1666464484
transform 1 0 76720 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_676
timestamp 1666464484
transform 1 0 77056 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_740
timestamp 1666464484
transform 1 0 84224 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_744
timestamp 1666464484
transform 1 0 84672 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_747
timestamp 1666464484
transform 1 0 85008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_811
timestamp 1666464484
transform 1 0 92176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_815
timestamp 1666464484
transform 1 0 92624 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_818
timestamp 1666464484
transform 1 0 92960 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_882
timestamp 1666464484
transform 1 0 100128 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_886
timestamp 1666464484
transform 1 0 100576 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_889
timestamp 1666464484
transform 1 0 100912 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_953
timestamp 1666464484
transform 1 0 108080 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_957
timestamp 1666464484
transform 1 0 108528 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_960
timestamp 1666464484
transform 1 0 108864 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1024
timestamp 1666464484
transform 1 0 116032 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1028
timestamp 1666464484
transform 1 0 116480 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_1031
timestamp 1666464484
transform 1 0 116816 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1095
timestamp 1666464484
transform 1 0 123984 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1099
timestamp 1666464484
transform 1 0 124432 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_1102
timestamp 1666464484
transform 1 0 124768 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1166
timestamp 1666464484
transform 1 0 131936 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1170
timestamp 1666464484
transform 1 0 132384 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_1173
timestamp 1666464484
transform 1 0 132720 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1237
timestamp 1666464484
transform 1 0 139888 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1241
timestamp 1666464484
transform 1 0 140336 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_1244
timestamp 1666464484
transform 1 0 140672 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1308
timestamp 1666464484
transform 1 0 147840 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1312
timestamp 1666464484
transform 1 0 148288 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_1315
timestamp 1666464484
transform 1 0 148624 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1379
timestamp 1666464484
transform 1 0 155792 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1383
timestamp 1666464484
transform 1 0 156240 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_1386
timestamp 1666464484
transform 1 0 156576 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1450
timestamp 1666464484
transform 1 0 163744 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1454
timestamp 1666464484
transform 1 0 164192 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_1457
timestamp 1666464484
transform 1 0 164528 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1521
timestamp 1666464484
transform 1 0 171696 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1525
timestamp 1666464484
transform 1 0 172144 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_1528
timestamp 1666464484
transform 1 0 172480 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_1560
timestamp 1666464484
transform 1 0 176064 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1576
timestamp 1666464484
transform 1 0 177856 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1580
timestamp 1666464484
transform 1 0 178304 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_2
timestamp 1666464484
transform 1 0 1568 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_66
timestamp 1666464484
transform 1 0 8736 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_70
timestamp 1666464484
transform 1 0 9184 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_73
timestamp 1666464484
transform 1 0 9520 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_137
timestamp 1666464484
transform 1 0 16688 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_141
timestamp 1666464484
transform 1 0 17136 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_144
timestamp 1666464484
transform 1 0 17472 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_208
timestamp 1666464484
transform 1 0 24640 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1666464484
transform 1 0 25088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_215
timestamp 1666464484
transform 1 0 25424 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_279
timestamp 1666464484
transform 1 0 32592 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1666464484
transform 1 0 33040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1666464484
transform 1 0 33376 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_350
timestamp 1666464484
transform 1 0 40544 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1666464484
transform 1 0 40992 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_357
timestamp 1666464484
transform 1 0 41328 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_421
timestamp 1666464484
transform 1 0 48496 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_425
timestamp 1666464484
transform 1 0 48944 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_428
timestamp 1666464484
transform 1 0 49280 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_492
timestamp 1666464484
transform 1 0 56448 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_496
timestamp 1666464484
transform 1 0 56896 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_499
timestamp 1666464484
transform 1 0 57232 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_563
timestamp 1666464484
transform 1 0 64400 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_567
timestamp 1666464484
transform 1 0 64848 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_570
timestamp 1666464484
transform 1 0 65184 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_634
timestamp 1666464484
transform 1 0 72352 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_638
timestamp 1666464484
transform 1 0 72800 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_641
timestamp 1666464484
transform 1 0 73136 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_705
timestamp 1666464484
transform 1 0 80304 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_709
timestamp 1666464484
transform 1 0 80752 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_712
timestamp 1666464484
transform 1 0 81088 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_776
timestamp 1666464484
transform 1 0 88256 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_780
timestamp 1666464484
transform 1 0 88704 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_783
timestamp 1666464484
transform 1 0 89040 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_847
timestamp 1666464484
transform 1 0 96208 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_851
timestamp 1666464484
transform 1 0 96656 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_854
timestamp 1666464484
transform 1 0 96992 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_918
timestamp 1666464484
transform 1 0 104160 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_922
timestamp 1666464484
transform 1 0 104608 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_925
timestamp 1666464484
transform 1 0 104944 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_989
timestamp 1666464484
transform 1 0 112112 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_993
timestamp 1666464484
transform 1 0 112560 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_996
timestamp 1666464484
transform 1 0 112896 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_1060
timestamp 1666464484
transform 1 0 120064 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1064
timestamp 1666464484
transform 1 0 120512 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_1067
timestamp 1666464484
transform 1 0 120848 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_1131
timestamp 1666464484
transform 1 0 128016 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1135
timestamp 1666464484
transform 1 0 128464 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_1138
timestamp 1666464484
transform 1 0 128800 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_1202
timestamp 1666464484
transform 1 0 135968 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1206
timestamp 1666464484
transform 1 0 136416 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_1209
timestamp 1666464484
transform 1 0 136752 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_1273
timestamp 1666464484
transform 1 0 143920 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1277
timestamp 1666464484
transform 1 0 144368 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_1280
timestamp 1666464484
transform 1 0 144704 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_1344
timestamp 1666464484
transform 1 0 151872 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1348
timestamp 1666464484
transform 1 0 152320 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_1351
timestamp 1666464484
transform 1 0 152656 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_1415
timestamp 1666464484
transform 1 0 159824 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1419
timestamp 1666464484
transform 1 0 160272 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_1422
timestamp 1666464484
transform 1 0 160608 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_1486
timestamp 1666464484
transform 1 0 167776 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1490
timestamp 1666464484
transform 1 0 168224 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_1493
timestamp 1666464484
transform 1 0 168560 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_1557
timestamp 1666464484
transform 1 0 175728 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1561
timestamp 1666464484
transform 1 0 176176 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_1564
timestamp 1666464484
transform 1 0 176512 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1580
timestamp 1666464484
transform 1 0 178304 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_2
timestamp 1666464484
transform 1 0 1568 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_34
timestamp 1666464484
transform 1 0 5152 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_37
timestamp 1666464484
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_101
timestamp 1666464484
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1666464484
transform 1 0 13104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_108
timestamp 1666464484
transform 1 0 13440 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_172
timestamp 1666464484
transform 1 0 20608 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1666464484
transform 1 0 21056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_179
timestamp 1666464484
transform 1 0 21392 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_243
timestamp 1666464484
transform 1 0 28560 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1666464484
transform 1 0 29008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_250
timestamp 1666464484
transform 1 0 29344 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_314
timestamp 1666464484
transform 1 0 36512 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_318
timestamp 1666464484
transform 1 0 36960 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1666464484
transform 1 0 37296 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_385
timestamp 1666464484
transform 1 0 44464 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1666464484
transform 1 0 44912 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_392
timestamp 1666464484
transform 1 0 45248 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_456
timestamp 1666464484
transform 1 0 52416 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_460
timestamp 1666464484
transform 1 0 52864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_463
timestamp 1666464484
transform 1 0 53200 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_527
timestamp 1666464484
transform 1 0 60368 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_531
timestamp 1666464484
transform 1 0 60816 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_534
timestamp 1666464484
transform 1 0 61152 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_598
timestamp 1666464484
transform 1 0 68320 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_602
timestamp 1666464484
transform 1 0 68768 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_605
timestamp 1666464484
transform 1 0 69104 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_669
timestamp 1666464484
transform 1 0 76272 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_673
timestamp 1666464484
transform 1 0 76720 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_676
timestamp 1666464484
transform 1 0 77056 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_740
timestamp 1666464484
transform 1 0 84224 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_744
timestamp 1666464484
transform 1 0 84672 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_747
timestamp 1666464484
transform 1 0 85008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_811
timestamp 1666464484
transform 1 0 92176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_815
timestamp 1666464484
transform 1 0 92624 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_818
timestamp 1666464484
transform 1 0 92960 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_882
timestamp 1666464484
transform 1 0 100128 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_886
timestamp 1666464484
transform 1 0 100576 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_889
timestamp 1666464484
transform 1 0 100912 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_953
timestamp 1666464484
transform 1 0 108080 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_957
timestamp 1666464484
transform 1 0 108528 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_960
timestamp 1666464484
transform 1 0 108864 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1024
timestamp 1666464484
transform 1 0 116032 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1028
timestamp 1666464484
transform 1 0 116480 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_1031
timestamp 1666464484
transform 1 0 116816 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1095
timestamp 1666464484
transform 1 0 123984 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1099
timestamp 1666464484
transform 1 0 124432 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_1102
timestamp 1666464484
transform 1 0 124768 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1166
timestamp 1666464484
transform 1 0 131936 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1170
timestamp 1666464484
transform 1 0 132384 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_1173
timestamp 1666464484
transform 1 0 132720 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1237
timestamp 1666464484
transform 1 0 139888 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1241
timestamp 1666464484
transform 1 0 140336 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_1244
timestamp 1666464484
transform 1 0 140672 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1308
timestamp 1666464484
transform 1 0 147840 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1312
timestamp 1666464484
transform 1 0 148288 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_1315
timestamp 1666464484
transform 1 0 148624 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1379
timestamp 1666464484
transform 1 0 155792 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1383
timestamp 1666464484
transform 1 0 156240 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_1386
timestamp 1666464484
transform 1 0 156576 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1450
timestamp 1666464484
transform 1 0 163744 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1454
timestamp 1666464484
transform 1 0 164192 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_1457
timestamp 1666464484
transform 1 0 164528 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1521
timestamp 1666464484
transform 1 0 171696 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1525
timestamp 1666464484
transform 1 0 172144 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_1528
timestamp 1666464484
transform 1 0 172480 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_1560
timestamp 1666464484
transform 1 0 176064 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1576
timestamp 1666464484
transform 1 0 177856 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1580
timestamp 1666464484
transform 1 0 178304 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_2
timestamp 1666464484
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_66
timestamp 1666464484
transform 1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_70
timestamp 1666464484
transform 1 0 9184 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_73
timestamp 1666464484
transform 1 0 9520 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_137
timestamp 1666464484
transform 1 0 16688 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1666464484
transform 1 0 17136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_144
timestamp 1666464484
transform 1 0 17472 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_208
timestamp 1666464484
transform 1 0 24640 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1666464484
transform 1 0 25088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_215
timestamp 1666464484
transform 1 0 25424 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_279
timestamp 1666464484
transform 1 0 32592 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_283
timestamp 1666464484
transform 1 0 33040 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1666464484
transform 1 0 33376 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_350
timestamp 1666464484
transform 1 0 40544 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1666464484
transform 1 0 40992 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_357
timestamp 1666464484
transform 1 0 41328 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_421
timestamp 1666464484
transform 1 0 48496 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_425
timestamp 1666464484
transform 1 0 48944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_428
timestamp 1666464484
transform 1 0 49280 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_492
timestamp 1666464484
transform 1 0 56448 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_496
timestamp 1666464484
transform 1 0 56896 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_499
timestamp 1666464484
transform 1 0 57232 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_563
timestamp 1666464484
transform 1 0 64400 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_567
timestamp 1666464484
transform 1 0 64848 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_570
timestamp 1666464484
transform 1 0 65184 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_634
timestamp 1666464484
transform 1 0 72352 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_638
timestamp 1666464484
transform 1 0 72800 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_641
timestamp 1666464484
transform 1 0 73136 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_705
timestamp 1666464484
transform 1 0 80304 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_709
timestamp 1666464484
transform 1 0 80752 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_712
timestamp 1666464484
transform 1 0 81088 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_776
timestamp 1666464484
transform 1 0 88256 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_780
timestamp 1666464484
transform 1 0 88704 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_783
timestamp 1666464484
transform 1 0 89040 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_847
timestamp 1666464484
transform 1 0 96208 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_851
timestamp 1666464484
transform 1 0 96656 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_854
timestamp 1666464484
transform 1 0 96992 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_918
timestamp 1666464484
transform 1 0 104160 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_922
timestamp 1666464484
transform 1 0 104608 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_925
timestamp 1666464484
transform 1 0 104944 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_989
timestamp 1666464484
transform 1 0 112112 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_993
timestamp 1666464484
transform 1 0 112560 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_996
timestamp 1666464484
transform 1 0 112896 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_1060
timestamp 1666464484
transform 1 0 120064 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1064
timestamp 1666464484
transform 1 0 120512 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_1067
timestamp 1666464484
transform 1 0 120848 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_1131
timestamp 1666464484
transform 1 0 128016 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1135
timestamp 1666464484
transform 1 0 128464 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_1138
timestamp 1666464484
transform 1 0 128800 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_1202
timestamp 1666464484
transform 1 0 135968 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1206
timestamp 1666464484
transform 1 0 136416 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_1209
timestamp 1666464484
transform 1 0 136752 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_1273
timestamp 1666464484
transform 1 0 143920 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1277
timestamp 1666464484
transform 1 0 144368 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_1280
timestamp 1666464484
transform 1 0 144704 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_1344
timestamp 1666464484
transform 1 0 151872 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1348
timestamp 1666464484
transform 1 0 152320 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_1351
timestamp 1666464484
transform 1 0 152656 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_1415
timestamp 1666464484
transform 1 0 159824 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1419
timestamp 1666464484
transform 1 0 160272 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_1422
timestamp 1666464484
transform 1 0 160608 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_1486
timestamp 1666464484
transform 1 0 167776 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1490
timestamp 1666464484
transform 1 0 168224 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_1493
timestamp 1666464484
transform 1 0 168560 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_1557
timestamp 1666464484
transform 1 0 175728 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1561
timestamp 1666464484
transform 1 0 176176 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_1564
timestamp 1666464484
transform 1 0 176512 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1580
timestamp 1666464484
transform 1 0 178304 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_2
timestamp 1666464484
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_34
timestamp 1666464484
transform 1 0 5152 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_37
timestamp 1666464484
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_101
timestamp 1666464484
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_105
timestamp 1666464484
transform 1 0 13104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_108
timestamp 1666464484
transform 1 0 13440 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_172
timestamp 1666464484
transform 1 0 20608 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_176
timestamp 1666464484
transform 1 0 21056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_179
timestamp 1666464484
transform 1 0 21392 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_243
timestamp 1666464484
transform 1 0 28560 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_247
timestamp 1666464484
transform 1 0 29008 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_250
timestamp 1666464484
transform 1 0 29344 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_314
timestamp 1666464484
transform 1 0 36512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1666464484
transform 1 0 36960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1666464484
transform 1 0 37296 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_385
timestamp 1666464484
transform 1 0 44464 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1666464484
transform 1 0 44912 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_392
timestamp 1666464484
transform 1 0 45248 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_456
timestamp 1666464484
transform 1 0 52416 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_460
timestamp 1666464484
transform 1 0 52864 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_463
timestamp 1666464484
transform 1 0 53200 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_527
timestamp 1666464484
transform 1 0 60368 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 60816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_534
timestamp 1666464484
transform 1 0 61152 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_598
timestamp 1666464484
transform 1 0 68320 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_602
timestamp 1666464484
transform 1 0 68768 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_605
timestamp 1666464484
transform 1 0 69104 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_669
timestamp 1666464484
transform 1 0 76272 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_673
timestamp 1666464484
transform 1 0 76720 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_676
timestamp 1666464484
transform 1 0 77056 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_740
timestamp 1666464484
transform 1 0 84224 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_744
timestamp 1666464484
transform 1 0 84672 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_747
timestamp 1666464484
transform 1 0 85008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_811
timestamp 1666464484
transform 1 0 92176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_815
timestamp 1666464484
transform 1 0 92624 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_818
timestamp 1666464484
transform 1 0 92960 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_882
timestamp 1666464484
transform 1 0 100128 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_886
timestamp 1666464484
transform 1 0 100576 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_889
timestamp 1666464484
transform 1 0 100912 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_953
timestamp 1666464484
transform 1 0 108080 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_957
timestamp 1666464484
transform 1 0 108528 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_960
timestamp 1666464484
transform 1 0 108864 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1024
timestamp 1666464484
transform 1 0 116032 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1028
timestamp 1666464484
transform 1 0 116480 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_1031
timestamp 1666464484
transform 1 0 116816 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1095
timestamp 1666464484
transform 1 0 123984 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1099
timestamp 1666464484
transform 1 0 124432 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_1102
timestamp 1666464484
transform 1 0 124768 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1166
timestamp 1666464484
transform 1 0 131936 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1170
timestamp 1666464484
transform 1 0 132384 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_1173
timestamp 1666464484
transform 1 0 132720 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1237
timestamp 1666464484
transform 1 0 139888 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1241
timestamp 1666464484
transform 1 0 140336 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_1244
timestamp 1666464484
transform 1 0 140672 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1308
timestamp 1666464484
transform 1 0 147840 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1312
timestamp 1666464484
transform 1 0 148288 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_1315
timestamp 1666464484
transform 1 0 148624 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1379
timestamp 1666464484
transform 1 0 155792 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1383
timestamp 1666464484
transform 1 0 156240 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_1386
timestamp 1666464484
transform 1 0 156576 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1450
timestamp 1666464484
transform 1 0 163744 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1454
timestamp 1666464484
transform 1 0 164192 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_1457
timestamp 1666464484
transform 1 0 164528 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1521
timestamp 1666464484
transform 1 0 171696 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1525
timestamp 1666464484
transform 1 0 172144 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_1528
timestamp 1666464484
transform 1 0 172480 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_1560
timestamp 1666464484
transform 1 0 176064 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1576
timestamp 1666464484
transform 1 0 177856 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1580
timestamp 1666464484
transform 1 0 178304 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_2
timestamp 1666464484
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_66
timestamp 1666464484
transform 1 0 8736 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_70
timestamp 1666464484
transform 1 0 9184 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_73
timestamp 1666464484
transform 1 0 9520 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_137
timestamp 1666464484
transform 1 0 16688 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_141
timestamp 1666464484
transform 1 0 17136 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_144
timestamp 1666464484
transform 1 0 17472 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_208
timestamp 1666464484
transform 1 0 24640 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1666464484
transform 1 0 25088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_215
timestamp 1666464484
transform 1 0 25424 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_279
timestamp 1666464484
transform 1 0 32592 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1666464484
transform 1 0 33040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1666464484
transform 1 0 33376 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_350
timestamp 1666464484
transform 1 0 40544 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1666464484
transform 1 0 40992 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_357
timestamp 1666464484
transform 1 0 41328 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_421
timestamp 1666464484
transform 1 0 48496 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_425
timestamp 1666464484
transform 1 0 48944 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_428
timestamp 1666464484
transform 1 0 49280 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_492
timestamp 1666464484
transform 1 0 56448 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_496
timestamp 1666464484
transform 1 0 56896 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_499
timestamp 1666464484
transform 1 0 57232 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_563
timestamp 1666464484
transform 1 0 64400 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_567
timestamp 1666464484
transform 1 0 64848 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_570
timestamp 1666464484
transform 1 0 65184 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_634
timestamp 1666464484
transform 1 0 72352 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_638
timestamp 1666464484
transform 1 0 72800 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_641
timestamp 1666464484
transform 1 0 73136 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_705
timestamp 1666464484
transform 1 0 80304 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_709
timestamp 1666464484
transform 1 0 80752 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_712
timestamp 1666464484
transform 1 0 81088 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_776
timestamp 1666464484
transform 1 0 88256 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_780
timestamp 1666464484
transform 1 0 88704 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_783
timestamp 1666464484
transform 1 0 89040 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_847
timestamp 1666464484
transform 1 0 96208 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_851
timestamp 1666464484
transform 1 0 96656 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_854
timestamp 1666464484
transform 1 0 96992 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_918
timestamp 1666464484
transform 1 0 104160 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_922
timestamp 1666464484
transform 1 0 104608 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_925
timestamp 1666464484
transform 1 0 104944 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_989
timestamp 1666464484
transform 1 0 112112 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_993
timestamp 1666464484
transform 1 0 112560 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_996
timestamp 1666464484
transform 1 0 112896 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_1060
timestamp 1666464484
transform 1 0 120064 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1064
timestamp 1666464484
transform 1 0 120512 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_1067
timestamp 1666464484
transform 1 0 120848 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_1131
timestamp 1666464484
transform 1 0 128016 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1135
timestamp 1666464484
transform 1 0 128464 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_1138
timestamp 1666464484
transform 1 0 128800 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_1202
timestamp 1666464484
transform 1 0 135968 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1206
timestamp 1666464484
transform 1 0 136416 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_1209
timestamp 1666464484
transform 1 0 136752 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_1273
timestamp 1666464484
transform 1 0 143920 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1277
timestamp 1666464484
transform 1 0 144368 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_1280
timestamp 1666464484
transform 1 0 144704 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_1344
timestamp 1666464484
transform 1 0 151872 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1348
timestamp 1666464484
transform 1 0 152320 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_1351
timestamp 1666464484
transform 1 0 152656 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_1415
timestamp 1666464484
transform 1 0 159824 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1419
timestamp 1666464484
transform 1 0 160272 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_1422
timestamp 1666464484
transform 1 0 160608 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_1486
timestamp 1666464484
transform 1 0 167776 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1490
timestamp 1666464484
transform 1 0 168224 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_1493
timestamp 1666464484
transform 1 0 168560 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_1557
timestamp 1666464484
transform 1 0 175728 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1561
timestamp 1666464484
transform 1 0 176176 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_1564
timestamp 1666464484
transform 1 0 176512 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1580
timestamp 1666464484
transform 1 0 178304 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_2
timestamp 1666464484
transform 1 0 1568 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_34
timestamp 1666464484
transform 1 0 5152 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_37
timestamp 1666464484
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_101
timestamp 1666464484
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_105
timestamp 1666464484
transform 1 0 13104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_108
timestamp 1666464484
transform 1 0 13440 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_172
timestamp 1666464484
transform 1 0 20608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_176
timestamp 1666464484
transform 1 0 21056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_179
timestamp 1666464484
transform 1 0 21392 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_243
timestamp 1666464484
transform 1 0 28560 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_247
timestamp 1666464484
transform 1 0 29008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_250
timestamp 1666464484
transform 1 0 29344 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_314
timestamp 1666464484
transform 1 0 36512 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_318
timestamp 1666464484
transform 1 0 36960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_321
timestamp 1666464484
transform 1 0 37296 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_385
timestamp 1666464484
transform 1 0 44464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_389
timestamp 1666464484
transform 1 0 44912 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_392
timestamp 1666464484
transform 1 0 45248 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_456
timestamp 1666464484
transform 1 0 52416 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_460
timestamp 1666464484
transform 1 0 52864 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_463
timestamp 1666464484
transform 1 0 53200 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_527
timestamp 1666464484
transform 1 0 60368 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 60816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_534
timestamp 1666464484
transform 1 0 61152 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_598
timestamp 1666464484
transform 1 0 68320 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_602
timestamp 1666464484
transform 1 0 68768 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_605
timestamp 1666464484
transform 1 0 69104 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_669
timestamp 1666464484
transform 1 0 76272 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_673
timestamp 1666464484
transform 1 0 76720 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_676
timestamp 1666464484
transform 1 0 77056 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_740
timestamp 1666464484
transform 1 0 84224 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_744
timestamp 1666464484
transform 1 0 84672 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_747
timestamp 1666464484
transform 1 0 85008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_811
timestamp 1666464484
transform 1 0 92176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_815
timestamp 1666464484
transform 1 0 92624 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_818
timestamp 1666464484
transform 1 0 92960 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_882
timestamp 1666464484
transform 1 0 100128 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_886
timestamp 1666464484
transform 1 0 100576 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_889
timestamp 1666464484
transform 1 0 100912 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_953
timestamp 1666464484
transform 1 0 108080 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_957
timestamp 1666464484
transform 1 0 108528 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_960
timestamp 1666464484
transform 1 0 108864 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1024
timestamp 1666464484
transform 1 0 116032 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1028
timestamp 1666464484
transform 1 0 116480 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_1031
timestamp 1666464484
transform 1 0 116816 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1095
timestamp 1666464484
transform 1 0 123984 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1099
timestamp 1666464484
transform 1 0 124432 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_1102
timestamp 1666464484
transform 1 0 124768 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1166
timestamp 1666464484
transform 1 0 131936 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1170
timestamp 1666464484
transform 1 0 132384 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_1173
timestamp 1666464484
transform 1 0 132720 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1237
timestamp 1666464484
transform 1 0 139888 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1241
timestamp 1666464484
transform 1 0 140336 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_1244
timestamp 1666464484
transform 1 0 140672 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1308
timestamp 1666464484
transform 1 0 147840 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1312
timestamp 1666464484
transform 1 0 148288 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_1315
timestamp 1666464484
transform 1 0 148624 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1379
timestamp 1666464484
transform 1 0 155792 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1383
timestamp 1666464484
transform 1 0 156240 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_1386
timestamp 1666464484
transform 1 0 156576 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1450
timestamp 1666464484
transform 1 0 163744 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1454
timestamp 1666464484
transform 1 0 164192 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_1457
timestamp 1666464484
transform 1 0 164528 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1521
timestamp 1666464484
transform 1 0 171696 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1525
timestamp 1666464484
transform 1 0 172144 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_1528
timestamp 1666464484
transform 1 0 172480 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_1560
timestamp 1666464484
transform 1 0 176064 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1576
timestamp 1666464484
transform 1 0 177856 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1580
timestamp 1666464484
transform 1 0 178304 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_2
timestamp 1666464484
transform 1 0 1568 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_66
timestamp 1666464484
transform 1 0 8736 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_70
timestamp 1666464484
transform 1 0 9184 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_73
timestamp 1666464484
transform 1 0 9520 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_137
timestamp 1666464484
transform 1 0 16688 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_141
timestamp 1666464484
transform 1 0 17136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_144
timestamp 1666464484
transform 1 0 17472 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_208
timestamp 1666464484
transform 1 0 24640 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_212
timestamp 1666464484
transform 1 0 25088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_215
timestamp 1666464484
transform 1 0 25424 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_279
timestamp 1666464484
transform 1 0 32592 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_283
timestamp 1666464484
transform 1 0 33040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_286
timestamp 1666464484
transform 1 0 33376 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_350
timestamp 1666464484
transform 1 0 40544 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_354
timestamp 1666464484
transform 1 0 40992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_357
timestamp 1666464484
transform 1 0 41328 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_421
timestamp 1666464484
transform 1 0 48496 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_425
timestamp 1666464484
transform 1 0 48944 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_428
timestamp 1666464484
transform 1 0 49280 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_492
timestamp 1666464484
transform 1 0 56448 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_496
timestamp 1666464484
transform 1 0 56896 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_499
timestamp 1666464484
transform 1 0 57232 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_563
timestamp 1666464484
transform 1 0 64400 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_567
timestamp 1666464484
transform 1 0 64848 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_570
timestamp 1666464484
transform 1 0 65184 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_634
timestamp 1666464484
transform 1 0 72352 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_638
timestamp 1666464484
transform 1 0 72800 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_641
timestamp 1666464484
transform 1 0 73136 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_705
timestamp 1666464484
transform 1 0 80304 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_709
timestamp 1666464484
transform 1 0 80752 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_712
timestamp 1666464484
transform 1 0 81088 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_776
timestamp 1666464484
transform 1 0 88256 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_780
timestamp 1666464484
transform 1 0 88704 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_783
timestamp 1666464484
transform 1 0 89040 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_847
timestamp 1666464484
transform 1 0 96208 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_851
timestamp 1666464484
transform 1 0 96656 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_854
timestamp 1666464484
transform 1 0 96992 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_918
timestamp 1666464484
transform 1 0 104160 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_922
timestamp 1666464484
transform 1 0 104608 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_925
timestamp 1666464484
transform 1 0 104944 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_989
timestamp 1666464484
transform 1 0 112112 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_993
timestamp 1666464484
transform 1 0 112560 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_996
timestamp 1666464484
transform 1 0 112896 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1060
timestamp 1666464484
transform 1 0 120064 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1064
timestamp 1666464484
transform 1 0 120512 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_1067
timestamp 1666464484
transform 1 0 120848 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1131
timestamp 1666464484
transform 1 0 128016 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1135
timestamp 1666464484
transform 1 0 128464 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_1138
timestamp 1666464484
transform 1 0 128800 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1202
timestamp 1666464484
transform 1 0 135968 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1206
timestamp 1666464484
transform 1 0 136416 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_1209
timestamp 1666464484
transform 1 0 136752 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1273
timestamp 1666464484
transform 1 0 143920 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1277
timestamp 1666464484
transform 1 0 144368 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_1280
timestamp 1666464484
transform 1 0 144704 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1344
timestamp 1666464484
transform 1 0 151872 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1348
timestamp 1666464484
transform 1 0 152320 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_1351
timestamp 1666464484
transform 1 0 152656 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1415
timestamp 1666464484
transform 1 0 159824 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1419
timestamp 1666464484
transform 1 0 160272 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_1422
timestamp 1666464484
transform 1 0 160608 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1486
timestamp 1666464484
transform 1 0 167776 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1490
timestamp 1666464484
transform 1 0 168224 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_1493
timestamp 1666464484
transform 1 0 168560 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_1557
timestamp 1666464484
transform 1 0 175728 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1561
timestamp 1666464484
transform 1 0 176176 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_1564
timestamp 1666464484
transform 1 0 176512 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1580
timestamp 1666464484
transform 1 0 178304 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_2
timestamp 1666464484
transform 1 0 1568 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_34
timestamp 1666464484
transform 1 0 5152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_37
timestamp 1666464484
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_101
timestamp 1666464484
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_105
timestamp 1666464484
transform 1 0 13104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_108
timestamp 1666464484
transform 1 0 13440 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_172
timestamp 1666464484
transform 1 0 20608 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_176
timestamp 1666464484
transform 1 0 21056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_179
timestamp 1666464484
transform 1 0 21392 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_243
timestamp 1666464484
transform 1 0 28560 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_247
timestamp 1666464484
transform 1 0 29008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_250
timestamp 1666464484
transform 1 0 29344 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_314
timestamp 1666464484
transform 1 0 36512 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_318
timestamp 1666464484
transform 1 0 36960 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_321
timestamp 1666464484
transform 1 0 37296 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_385
timestamp 1666464484
transform 1 0 44464 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_389
timestamp 1666464484
transform 1 0 44912 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_392
timestamp 1666464484
transform 1 0 45248 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_456
timestamp 1666464484
transform 1 0 52416 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_460
timestamp 1666464484
transform 1 0 52864 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_463
timestamp 1666464484
transform 1 0 53200 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_527
timestamp 1666464484
transform 1 0 60368 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_531
timestamp 1666464484
transform 1 0 60816 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_534
timestamp 1666464484
transform 1 0 61152 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_598
timestamp 1666464484
transform 1 0 68320 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_602
timestamp 1666464484
transform 1 0 68768 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_605
timestamp 1666464484
transform 1 0 69104 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_669
timestamp 1666464484
transform 1 0 76272 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_673
timestamp 1666464484
transform 1 0 76720 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_676
timestamp 1666464484
transform 1 0 77056 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_740
timestamp 1666464484
transform 1 0 84224 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_744
timestamp 1666464484
transform 1 0 84672 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_747
timestamp 1666464484
transform 1 0 85008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_811
timestamp 1666464484
transform 1 0 92176 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_815
timestamp 1666464484
transform 1 0 92624 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_818
timestamp 1666464484
transform 1 0 92960 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_882
timestamp 1666464484
transform 1 0 100128 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_886
timestamp 1666464484
transform 1 0 100576 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_889
timestamp 1666464484
transform 1 0 100912 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_953
timestamp 1666464484
transform 1 0 108080 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_957
timestamp 1666464484
transform 1 0 108528 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_960
timestamp 1666464484
transform 1 0 108864 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1024
timestamp 1666464484
transform 1 0 116032 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1028
timestamp 1666464484
transform 1 0 116480 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_1031
timestamp 1666464484
transform 1 0 116816 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1095
timestamp 1666464484
transform 1 0 123984 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1099
timestamp 1666464484
transform 1 0 124432 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_1102
timestamp 1666464484
transform 1 0 124768 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1166
timestamp 1666464484
transform 1 0 131936 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1170
timestamp 1666464484
transform 1 0 132384 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_1173
timestamp 1666464484
transform 1 0 132720 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1237
timestamp 1666464484
transform 1 0 139888 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1241
timestamp 1666464484
transform 1 0 140336 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_1244
timestamp 1666464484
transform 1 0 140672 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1308
timestamp 1666464484
transform 1 0 147840 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1312
timestamp 1666464484
transform 1 0 148288 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_1315
timestamp 1666464484
transform 1 0 148624 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1379
timestamp 1666464484
transform 1 0 155792 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1383
timestamp 1666464484
transform 1 0 156240 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_1386
timestamp 1666464484
transform 1 0 156576 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1450
timestamp 1666464484
transform 1 0 163744 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1454
timestamp 1666464484
transform 1 0 164192 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_1457
timestamp 1666464484
transform 1 0 164528 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1521
timestamp 1666464484
transform 1 0 171696 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1525
timestamp 1666464484
transform 1 0 172144 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_1528
timestamp 1666464484
transform 1 0 172480 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_1560
timestamp 1666464484
transform 1 0 176064 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1576
timestamp 1666464484
transform 1 0 177856 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1580
timestamp 1666464484
transform 1 0 178304 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_2
timestamp 1666464484
transform 1 0 1568 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_66
timestamp 1666464484
transform 1 0 8736 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_70
timestamp 1666464484
transform 1 0 9184 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_73
timestamp 1666464484
transform 1 0 9520 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_137
timestamp 1666464484
transform 1 0 16688 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_141
timestamp 1666464484
transform 1 0 17136 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_144
timestamp 1666464484
transform 1 0 17472 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_208
timestamp 1666464484
transform 1 0 24640 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_212
timestamp 1666464484
transform 1 0 25088 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_215
timestamp 1666464484
transform 1 0 25424 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_279
timestamp 1666464484
transform 1 0 32592 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_283
timestamp 1666464484
transform 1 0 33040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_286
timestamp 1666464484
transform 1 0 33376 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_350
timestamp 1666464484
transform 1 0 40544 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_354
timestamp 1666464484
transform 1 0 40992 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_357
timestamp 1666464484
transform 1 0 41328 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_421
timestamp 1666464484
transform 1 0 48496 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_425
timestamp 1666464484
transform 1 0 48944 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_428
timestamp 1666464484
transform 1 0 49280 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_492
timestamp 1666464484
transform 1 0 56448 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_496
timestamp 1666464484
transform 1 0 56896 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_499
timestamp 1666464484
transform 1 0 57232 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_563
timestamp 1666464484
transform 1 0 64400 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_567
timestamp 1666464484
transform 1 0 64848 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_570
timestamp 1666464484
transform 1 0 65184 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_634
timestamp 1666464484
transform 1 0 72352 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_638
timestamp 1666464484
transform 1 0 72800 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_641
timestamp 1666464484
transform 1 0 73136 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_705
timestamp 1666464484
transform 1 0 80304 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_709
timestamp 1666464484
transform 1 0 80752 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_712
timestamp 1666464484
transform 1 0 81088 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_776
timestamp 1666464484
transform 1 0 88256 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_780
timestamp 1666464484
transform 1 0 88704 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_783
timestamp 1666464484
transform 1 0 89040 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_847
timestamp 1666464484
transform 1 0 96208 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_851
timestamp 1666464484
transform 1 0 96656 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_854
timestamp 1666464484
transform 1 0 96992 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_918
timestamp 1666464484
transform 1 0 104160 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_922
timestamp 1666464484
transform 1 0 104608 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_925
timestamp 1666464484
transform 1 0 104944 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_989
timestamp 1666464484
transform 1 0 112112 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_993
timestamp 1666464484
transform 1 0 112560 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_996
timestamp 1666464484
transform 1 0 112896 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1060
timestamp 1666464484
transform 1 0 120064 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1064
timestamp 1666464484
transform 1 0 120512 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_1067
timestamp 1666464484
transform 1 0 120848 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1131
timestamp 1666464484
transform 1 0 128016 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1135
timestamp 1666464484
transform 1 0 128464 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_1138
timestamp 1666464484
transform 1 0 128800 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1202
timestamp 1666464484
transform 1 0 135968 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1206
timestamp 1666464484
transform 1 0 136416 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_1209
timestamp 1666464484
transform 1 0 136752 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1273
timestamp 1666464484
transform 1 0 143920 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1277
timestamp 1666464484
transform 1 0 144368 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_1280
timestamp 1666464484
transform 1 0 144704 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1344
timestamp 1666464484
transform 1 0 151872 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1348
timestamp 1666464484
transform 1 0 152320 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_1351
timestamp 1666464484
transform 1 0 152656 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1415
timestamp 1666464484
transform 1 0 159824 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1419
timestamp 1666464484
transform 1 0 160272 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_1422
timestamp 1666464484
transform 1 0 160608 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1486
timestamp 1666464484
transform 1 0 167776 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1490
timestamp 1666464484
transform 1 0 168224 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_1493
timestamp 1666464484
transform 1 0 168560 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1557
timestamp 1666464484
transform 1 0 175728 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1561
timestamp 1666464484
transform 1 0 176176 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_1564
timestamp 1666464484
transform 1 0 176512 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1580
timestamp 1666464484
transform 1 0 178304 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_2
timestamp 1666464484
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_34
timestamp 1666464484
transform 1 0 5152 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_37
timestamp 1666464484
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_101
timestamp 1666464484
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_105
timestamp 1666464484
transform 1 0 13104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_108
timestamp 1666464484
transform 1 0 13440 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_172
timestamp 1666464484
transform 1 0 20608 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_176
timestamp 1666464484
transform 1 0 21056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_179
timestamp 1666464484
transform 1 0 21392 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_243
timestamp 1666464484
transform 1 0 28560 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_247
timestamp 1666464484
transform 1 0 29008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_250
timestamp 1666464484
transform 1 0 29344 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_314
timestamp 1666464484
transform 1 0 36512 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_318
timestamp 1666464484
transform 1 0 36960 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_321
timestamp 1666464484
transform 1 0 37296 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_385
timestamp 1666464484
transform 1 0 44464 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_389
timestamp 1666464484
transform 1 0 44912 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_392
timestamp 1666464484
transform 1 0 45248 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_456
timestamp 1666464484
transform 1 0 52416 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_460
timestamp 1666464484
transform 1 0 52864 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_463
timestamp 1666464484
transform 1 0 53200 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_527
timestamp 1666464484
transform 1 0 60368 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 60816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_534
timestamp 1666464484
transform 1 0 61152 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_598
timestamp 1666464484
transform 1 0 68320 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_602
timestamp 1666464484
transform 1 0 68768 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_605
timestamp 1666464484
transform 1 0 69104 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_669
timestamp 1666464484
transform 1 0 76272 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_673
timestamp 1666464484
transform 1 0 76720 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_676
timestamp 1666464484
transform 1 0 77056 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_740
timestamp 1666464484
transform 1 0 84224 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_744
timestamp 1666464484
transform 1 0 84672 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_747
timestamp 1666464484
transform 1 0 85008 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_811
timestamp 1666464484
transform 1 0 92176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_815
timestamp 1666464484
transform 1 0 92624 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_818
timestamp 1666464484
transform 1 0 92960 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_882
timestamp 1666464484
transform 1 0 100128 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_886
timestamp 1666464484
transform 1 0 100576 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_889
timestamp 1666464484
transform 1 0 100912 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_953
timestamp 1666464484
transform 1 0 108080 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_957
timestamp 1666464484
transform 1 0 108528 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_960
timestamp 1666464484
transform 1 0 108864 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1024
timestamp 1666464484
transform 1 0 116032 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1028
timestamp 1666464484
transform 1 0 116480 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_1031
timestamp 1666464484
transform 1 0 116816 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1095
timestamp 1666464484
transform 1 0 123984 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1099
timestamp 1666464484
transform 1 0 124432 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_1102
timestamp 1666464484
transform 1 0 124768 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1166
timestamp 1666464484
transform 1 0 131936 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1170
timestamp 1666464484
transform 1 0 132384 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_1173
timestamp 1666464484
transform 1 0 132720 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1237
timestamp 1666464484
transform 1 0 139888 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1241
timestamp 1666464484
transform 1 0 140336 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_1244
timestamp 1666464484
transform 1 0 140672 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1308
timestamp 1666464484
transform 1 0 147840 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1312
timestamp 1666464484
transform 1 0 148288 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_1315
timestamp 1666464484
transform 1 0 148624 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1379
timestamp 1666464484
transform 1 0 155792 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1383
timestamp 1666464484
transform 1 0 156240 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_1386
timestamp 1666464484
transform 1 0 156576 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1450
timestamp 1666464484
transform 1 0 163744 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1454
timestamp 1666464484
transform 1 0 164192 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_1457
timestamp 1666464484
transform 1 0 164528 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1521
timestamp 1666464484
transform 1 0 171696 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1525
timestamp 1666464484
transform 1 0 172144 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_1528
timestamp 1666464484
transform 1 0 172480 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_1560
timestamp 1666464484
transform 1 0 176064 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1576
timestamp 1666464484
transform 1 0 177856 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1580
timestamp 1666464484
transform 1 0 178304 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_2
timestamp 1666464484
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_66
timestamp 1666464484
transform 1 0 8736 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_70
timestamp 1666464484
transform 1 0 9184 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_73
timestamp 1666464484
transform 1 0 9520 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_137
timestamp 1666464484
transform 1 0 16688 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_141
timestamp 1666464484
transform 1 0 17136 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_144
timestamp 1666464484
transform 1 0 17472 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_208
timestamp 1666464484
transform 1 0 24640 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_212
timestamp 1666464484
transform 1 0 25088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_215
timestamp 1666464484
transform 1 0 25424 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_279
timestamp 1666464484
transform 1 0 32592 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_283
timestamp 1666464484
transform 1 0 33040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_286
timestamp 1666464484
transform 1 0 33376 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_350
timestamp 1666464484
transform 1 0 40544 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_354
timestamp 1666464484
transform 1 0 40992 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_357
timestamp 1666464484
transform 1 0 41328 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_421
timestamp 1666464484
transform 1 0 48496 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_425
timestamp 1666464484
transform 1 0 48944 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_428
timestamp 1666464484
transform 1 0 49280 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_492
timestamp 1666464484
transform 1 0 56448 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_496
timestamp 1666464484
transform 1 0 56896 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_499
timestamp 1666464484
transform 1 0 57232 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_563
timestamp 1666464484
transform 1 0 64400 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_567
timestamp 1666464484
transform 1 0 64848 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_570
timestamp 1666464484
transform 1 0 65184 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_634
timestamp 1666464484
transform 1 0 72352 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_638
timestamp 1666464484
transform 1 0 72800 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_641
timestamp 1666464484
transform 1 0 73136 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_705
timestamp 1666464484
transform 1 0 80304 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_709
timestamp 1666464484
transform 1 0 80752 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_712
timestamp 1666464484
transform 1 0 81088 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_776
timestamp 1666464484
transform 1 0 88256 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_780
timestamp 1666464484
transform 1 0 88704 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_783
timestamp 1666464484
transform 1 0 89040 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_847
timestamp 1666464484
transform 1 0 96208 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_851
timestamp 1666464484
transform 1 0 96656 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_854
timestamp 1666464484
transform 1 0 96992 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_918
timestamp 1666464484
transform 1 0 104160 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_922
timestamp 1666464484
transform 1 0 104608 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_925
timestamp 1666464484
transform 1 0 104944 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_989
timestamp 1666464484
transform 1 0 112112 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_993
timestamp 1666464484
transform 1 0 112560 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_996
timestamp 1666464484
transform 1 0 112896 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1060
timestamp 1666464484
transform 1 0 120064 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1064
timestamp 1666464484
transform 1 0 120512 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_1067
timestamp 1666464484
transform 1 0 120848 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1131
timestamp 1666464484
transform 1 0 128016 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1135
timestamp 1666464484
transform 1 0 128464 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_1138
timestamp 1666464484
transform 1 0 128800 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1202
timestamp 1666464484
transform 1 0 135968 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1206
timestamp 1666464484
transform 1 0 136416 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_1209
timestamp 1666464484
transform 1 0 136752 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1273
timestamp 1666464484
transform 1 0 143920 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1277
timestamp 1666464484
transform 1 0 144368 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_1280
timestamp 1666464484
transform 1 0 144704 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1344
timestamp 1666464484
transform 1 0 151872 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1348
timestamp 1666464484
transform 1 0 152320 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_1351
timestamp 1666464484
transform 1 0 152656 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1415
timestamp 1666464484
transform 1 0 159824 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1419
timestamp 1666464484
transform 1 0 160272 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_1422
timestamp 1666464484
transform 1 0 160608 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1486
timestamp 1666464484
transform 1 0 167776 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1490
timestamp 1666464484
transform 1 0 168224 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_1493
timestamp 1666464484
transform 1 0 168560 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_1557
timestamp 1666464484
transform 1 0 175728 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1561
timestamp 1666464484
transform 1 0 176176 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_1564
timestamp 1666464484
transform 1 0 176512 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1580
timestamp 1666464484
transform 1 0 178304 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_86_2
timestamp 1666464484
transform 1 0 1568 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_34
timestamp 1666464484
transform 1 0 5152 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_37
timestamp 1666464484
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_101
timestamp 1666464484
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_105
timestamp 1666464484
transform 1 0 13104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_108
timestamp 1666464484
transform 1 0 13440 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_172
timestamp 1666464484
transform 1 0 20608 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_176
timestamp 1666464484
transform 1 0 21056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_179
timestamp 1666464484
transform 1 0 21392 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_243
timestamp 1666464484
transform 1 0 28560 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_247
timestamp 1666464484
transform 1 0 29008 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_250
timestamp 1666464484
transform 1 0 29344 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_314
timestamp 1666464484
transform 1 0 36512 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_318
timestamp 1666464484
transform 1 0 36960 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_321
timestamp 1666464484
transform 1 0 37296 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_385
timestamp 1666464484
transform 1 0 44464 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_389
timestamp 1666464484
transform 1 0 44912 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_392
timestamp 1666464484
transform 1 0 45248 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_456
timestamp 1666464484
transform 1 0 52416 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_460
timestamp 1666464484
transform 1 0 52864 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_463
timestamp 1666464484
transform 1 0 53200 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_527
timestamp 1666464484
transform 1 0 60368 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 60816 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_534
timestamp 1666464484
transform 1 0 61152 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_598
timestamp 1666464484
transform 1 0 68320 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_602
timestamp 1666464484
transform 1 0 68768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_605
timestamp 1666464484
transform 1 0 69104 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_669
timestamp 1666464484
transform 1 0 76272 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_673
timestamp 1666464484
transform 1 0 76720 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_676
timestamp 1666464484
transform 1 0 77056 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_740
timestamp 1666464484
transform 1 0 84224 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_744
timestamp 1666464484
transform 1 0 84672 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_747
timestamp 1666464484
transform 1 0 85008 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_811
timestamp 1666464484
transform 1 0 92176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_815
timestamp 1666464484
transform 1 0 92624 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_818
timestamp 1666464484
transform 1 0 92960 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_882
timestamp 1666464484
transform 1 0 100128 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_886
timestamp 1666464484
transform 1 0 100576 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_889
timestamp 1666464484
transform 1 0 100912 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_953
timestamp 1666464484
transform 1 0 108080 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_957
timestamp 1666464484
transform 1 0 108528 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_960
timestamp 1666464484
transform 1 0 108864 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1024
timestamp 1666464484
transform 1 0 116032 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1028
timestamp 1666464484
transform 1 0 116480 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_1031
timestamp 1666464484
transform 1 0 116816 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1095
timestamp 1666464484
transform 1 0 123984 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1099
timestamp 1666464484
transform 1 0 124432 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_1102
timestamp 1666464484
transform 1 0 124768 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1166
timestamp 1666464484
transform 1 0 131936 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1170
timestamp 1666464484
transform 1 0 132384 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_1173
timestamp 1666464484
transform 1 0 132720 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1237
timestamp 1666464484
transform 1 0 139888 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1241
timestamp 1666464484
transform 1 0 140336 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_1244
timestamp 1666464484
transform 1 0 140672 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1308
timestamp 1666464484
transform 1 0 147840 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1312
timestamp 1666464484
transform 1 0 148288 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_1315
timestamp 1666464484
transform 1 0 148624 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1379
timestamp 1666464484
transform 1 0 155792 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1383
timestamp 1666464484
transform 1 0 156240 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_1386
timestamp 1666464484
transform 1 0 156576 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1450
timestamp 1666464484
transform 1 0 163744 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1454
timestamp 1666464484
transform 1 0 164192 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_1457
timestamp 1666464484
transform 1 0 164528 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1521
timestamp 1666464484
transform 1 0 171696 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1525
timestamp 1666464484
transform 1 0 172144 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_86_1528
timestamp 1666464484
transform 1 0 172480 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_1560
timestamp 1666464484
transform 1 0 176064 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1576
timestamp 1666464484
transform 1 0 177856 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1580
timestamp 1666464484
transform 1 0 178304 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_2
timestamp 1666464484
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_66
timestamp 1666464484
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_70
timestamp 1666464484
transform 1 0 9184 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_73
timestamp 1666464484
transform 1 0 9520 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_137
timestamp 1666464484
transform 1 0 16688 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_141
timestamp 1666464484
transform 1 0 17136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_144
timestamp 1666464484
transform 1 0 17472 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_208
timestamp 1666464484
transform 1 0 24640 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_212
timestamp 1666464484
transform 1 0 25088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_215
timestamp 1666464484
transform 1 0 25424 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_279
timestamp 1666464484
transform 1 0 32592 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_283
timestamp 1666464484
transform 1 0 33040 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_286
timestamp 1666464484
transform 1 0 33376 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_350
timestamp 1666464484
transform 1 0 40544 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_354
timestamp 1666464484
transform 1 0 40992 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_357
timestamp 1666464484
transform 1 0 41328 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_421
timestamp 1666464484
transform 1 0 48496 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_425
timestamp 1666464484
transform 1 0 48944 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_428
timestamp 1666464484
transform 1 0 49280 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_492
timestamp 1666464484
transform 1 0 56448 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_496
timestamp 1666464484
transform 1 0 56896 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_499
timestamp 1666464484
transform 1 0 57232 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_563
timestamp 1666464484
transform 1 0 64400 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_567
timestamp 1666464484
transform 1 0 64848 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_570
timestamp 1666464484
transform 1 0 65184 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_634
timestamp 1666464484
transform 1 0 72352 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_638
timestamp 1666464484
transform 1 0 72800 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_641
timestamp 1666464484
transform 1 0 73136 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_705
timestamp 1666464484
transform 1 0 80304 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_709
timestamp 1666464484
transform 1 0 80752 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_712
timestamp 1666464484
transform 1 0 81088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_776
timestamp 1666464484
transform 1 0 88256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_780
timestamp 1666464484
transform 1 0 88704 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_783
timestamp 1666464484
transform 1 0 89040 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_847
timestamp 1666464484
transform 1 0 96208 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_851
timestamp 1666464484
transform 1 0 96656 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_854
timestamp 1666464484
transform 1 0 96992 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_918
timestamp 1666464484
transform 1 0 104160 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_922
timestamp 1666464484
transform 1 0 104608 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_925
timestamp 1666464484
transform 1 0 104944 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_989
timestamp 1666464484
transform 1 0 112112 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_993
timestamp 1666464484
transform 1 0 112560 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_996
timestamp 1666464484
transform 1 0 112896 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_1060
timestamp 1666464484
transform 1 0 120064 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1064
timestamp 1666464484
transform 1 0 120512 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_1067
timestamp 1666464484
transform 1 0 120848 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_1131
timestamp 1666464484
transform 1 0 128016 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1135
timestamp 1666464484
transform 1 0 128464 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_1138
timestamp 1666464484
transform 1 0 128800 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_1202
timestamp 1666464484
transform 1 0 135968 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1206
timestamp 1666464484
transform 1 0 136416 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_1209
timestamp 1666464484
transform 1 0 136752 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_1273
timestamp 1666464484
transform 1 0 143920 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1277
timestamp 1666464484
transform 1 0 144368 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_1280
timestamp 1666464484
transform 1 0 144704 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_1344
timestamp 1666464484
transform 1 0 151872 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1348
timestamp 1666464484
transform 1 0 152320 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_1351
timestamp 1666464484
transform 1 0 152656 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_1415
timestamp 1666464484
transform 1 0 159824 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1419
timestamp 1666464484
transform 1 0 160272 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_1422
timestamp 1666464484
transform 1 0 160608 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_1486
timestamp 1666464484
transform 1 0 167776 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1490
timestamp 1666464484
transform 1 0 168224 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_1493
timestamp 1666464484
transform 1 0 168560 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_1557
timestamp 1666464484
transform 1 0 175728 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1561
timestamp 1666464484
transform 1 0 176176 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_1564
timestamp 1666464484
transform 1 0 176512 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1580
timestamp 1666464484
transform 1 0 178304 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_2
timestamp 1666464484
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_34
timestamp 1666464484
transform 1 0 5152 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_37
timestamp 1666464484
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_101
timestamp 1666464484
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_105
timestamp 1666464484
transform 1 0 13104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_108
timestamp 1666464484
transform 1 0 13440 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_172
timestamp 1666464484
transform 1 0 20608 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_176
timestamp 1666464484
transform 1 0 21056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_179
timestamp 1666464484
transform 1 0 21392 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_243
timestamp 1666464484
transform 1 0 28560 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_247
timestamp 1666464484
transform 1 0 29008 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_250
timestamp 1666464484
transform 1 0 29344 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_314
timestamp 1666464484
transform 1 0 36512 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_318
timestamp 1666464484
transform 1 0 36960 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_321
timestamp 1666464484
transform 1 0 37296 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_385
timestamp 1666464484
transform 1 0 44464 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_389
timestamp 1666464484
transform 1 0 44912 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_392
timestamp 1666464484
transform 1 0 45248 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_456
timestamp 1666464484
transform 1 0 52416 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_460
timestamp 1666464484
transform 1 0 52864 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_463
timestamp 1666464484
transform 1 0 53200 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_527
timestamp 1666464484
transform 1 0 60368 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 60816 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_534
timestamp 1666464484
transform 1 0 61152 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_598
timestamp 1666464484
transform 1 0 68320 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_602
timestamp 1666464484
transform 1 0 68768 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_605
timestamp 1666464484
transform 1 0 69104 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_669
timestamp 1666464484
transform 1 0 76272 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_673
timestamp 1666464484
transform 1 0 76720 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_676
timestamp 1666464484
transform 1 0 77056 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_740
timestamp 1666464484
transform 1 0 84224 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_744
timestamp 1666464484
transform 1 0 84672 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_747
timestamp 1666464484
transform 1 0 85008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_811
timestamp 1666464484
transform 1 0 92176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_815
timestamp 1666464484
transform 1 0 92624 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_818
timestamp 1666464484
transform 1 0 92960 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_882
timestamp 1666464484
transform 1 0 100128 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_886
timestamp 1666464484
transform 1 0 100576 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_889
timestamp 1666464484
transform 1 0 100912 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_953
timestamp 1666464484
transform 1 0 108080 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_957
timestamp 1666464484
transform 1 0 108528 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_960
timestamp 1666464484
transform 1 0 108864 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1024
timestamp 1666464484
transform 1 0 116032 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1028
timestamp 1666464484
transform 1 0 116480 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_1031
timestamp 1666464484
transform 1 0 116816 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1095
timestamp 1666464484
transform 1 0 123984 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1099
timestamp 1666464484
transform 1 0 124432 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_1102
timestamp 1666464484
transform 1 0 124768 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1166
timestamp 1666464484
transform 1 0 131936 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1170
timestamp 1666464484
transform 1 0 132384 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_1173
timestamp 1666464484
transform 1 0 132720 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1237
timestamp 1666464484
transform 1 0 139888 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1241
timestamp 1666464484
transform 1 0 140336 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_1244
timestamp 1666464484
transform 1 0 140672 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1308
timestamp 1666464484
transform 1 0 147840 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1312
timestamp 1666464484
transform 1 0 148288 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_1315
timestamp 1666464484
transform 1 0 148624 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1379
timestamp 1666464484
transform 1 0 155792 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1383
timestamp 1666464484
transform 1 0 156240 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_1386
timestamp 1666464484
transform 1 0 156576 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1450
timestamp 1666464484
transform 1 0 163744 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1454
timestamp 1666464484
transform 1 0 164192 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_1457
timestamp 1666464484
transform 1 0 164528 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1521
timestamp 1666464484
transform 1 0 171696 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1525
timestamp 1666464484
transform 1 0 172144 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_1528
timestamp 1666464484
transform 1 0 172480 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_1560
timestamp 1666464484
transform 1 0 176064 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1576
timestamp 1666464484
transform 1 0 177856 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1580
timestamp 1666464484
transform 1 0 178304 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_2
timestamp 1666464484
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_66
timestamp 1666464484
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_70
timestamp 1666464484
transform 1 0 9184 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_73
timestamp 1666464484
transform 1 0 9520 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_137
timestamp 1666464484
transform 1 0 16688 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_141
timestamp 1666464484
transform 1 0 17136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_144
timestamp 1666464484
transform 1 0 17472 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_208
timestamp 1666464484
transform 1 0 24640 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_212
timestamp 1666464484
transform 1 0 25088 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_215
timestamp 1666464484
transform 1 0 25424 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_279
timestamp 1666464484
transform 1 0 32592 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_283
timestamp 1666464484
transform 1 0 33040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_286
timestamp 1666464484
transform 1 0 33376 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_350
timestamp 1666464484
transform 1 0 40544 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_354
timestamp 1666464484
transform 1 0 40992 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_357
timestamp 1666464484
transform 1 0 41328 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_421
timestamp 1666464484
transform 1 0 48496 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_425
timestamp 1666464484
transform 1 0 48944 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_428
timestamp 1666464484
transform 1 0 49280 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_492
timestamp 1666464484
transform 1 0 56448 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_496
timestamp 1666464484
transform 1 0 56896 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_499
timestamp 1666464484
transform 1 0 57232 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_563
timestamp 1666464484
transform 1 0 64400 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_567
timestamp 1666464484
transform 1 0 64848 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_570
timestamp 1666464484
transform 1 0 65184 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_634
timestamp 1666464484
transform 1 0 72352 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_638
timestamp 1666464484
transform 1 0 72800 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_641
timestamp 1666464484
transform 1 0 73136 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_705
timestamp 1666464484
transform 1 0 80304 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_709
timestamp 1666464484
transform 1 0 80752 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_712
timestamp 1666464484
transform 1 0 81088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_776
timestamp 1666464484
transform 1 0 88256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_780
timestamp 1666464484
transform 1 0 88704 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_783
timestamp 1666464484
transform 1 0 89040 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_847
timestamp 1666464484
transform 1 0 96208 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_851
timestamp 1666464484
transform 1 0 96656 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_854
timestamp 1666464484
transform 1 0 96992 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_918
timestamp 1666464484
transform 1 0 104160 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_922
timestamp 1666464484
transform 1 0 104608 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_925
timestamp 1666464484
transform 1 0 104944 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_989
timestamp 1666464484
transform 1 0 112112 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_993
timestamp 1666464484
transform 1 0 112560 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_996
timestamp 1666464484
transform 1 0 112896 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_1060
timestamp 1666464484
transform 1 0 120064 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1064
timestamp 1666464484
transform 1 0 120512 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_1067
timestamp 1666464484
transform 1 0 120848 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_1131
timestamp 1666464484
transform 1 0 128016 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1135
timestamp 1666464484
transform 1 0 128464 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_1138
timestamp 1666464484
transform 1 0 128800 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_1202
timestamp 1666464484
transform 1 0 135968 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1206
timestamp 1666464484
transform 1 0 136416 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_1209
timestamp 1666464484
transform 1 0 136752 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_1273
timestamp 1666464484
transform 1 0 143920 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1277
timestamp 1666464484
transform 1 0 144368 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_1280
timestamp 1666464484
transform 1 0 144704 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_1344
timestamp 1666464484
transform 1 0 151872 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1348
timestamp 1666464484
transform 1 0 152320 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_1351
timestamp 1666464484
transform 1 0 152656 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_1415
timestamp 1666464484
transform 1 0 159824 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1419
timestamp 1666464484
transform 1 0 160272 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_1422
timestamp 1666464484
transform 1 0 160608 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_1486
timestamp 1666464484
transform 1 0 167776 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1490
timestamp 1666464484
transform 1 0 168224 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_1493
timestamp 1666464484
transform 1 0 168560 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_1557
timestamp 1666464484
transform 1 0 175728 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1561
timestamp 1666464484
transform 1 0 176176 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_1564
timestamp 1666464484
transform 1 0 176512 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1580
timestamp 1666464484
transform 1 0 178304 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_2
timestamp 1666464484
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_34
timestamp 1666464484
transform 1 0 5152 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_37
timestamp 1666464484
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_101
timestamp 1666464484
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_105
timestamp 1666464484
transform 1 0 13104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_108
timestamp 1666464484
transform 1 0 13440 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_172
timestamp 1666464484
transform 1 0 20608 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_176
timestamp 1666464484
transform 1 0 21056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_179
timestamp 1666464484
transform 1 0 21392 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_243
timestamp 1666464484
transform 1 0 28560 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_247
timestamp 1666464484
transform 1 0 29008 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_250
timestamp 1666464484
transform 1 0 29344 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_314
timestamp 1666464484
transform 1 0 36512 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_318
timestamp 1666464484
transform 1 0 36960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_321
timestamp 1666464484
transform 1 0 37296 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_385
timestamp 1666464484
transform 1 0 44464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_389
timestamp 1666464484
transform 1 0 44912 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_392
timestamp 1666464484
transform 1 0 45248 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_456
timestamp 1666464484
transform 1 0 52416 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_460
timestamp 1666464484
transform 1 0 52864 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_463
timestamp 1666464484
transform 1 0 53200 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_527
timestamp 1666464484
transform 1 0 60368 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 60816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_534
timestamp 1666464484
transform 1 0 61152 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_598
timestamp 1666464484
transform 1 0 68320 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_602
timestamp 1666464484
transform 1 0 68768 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_605
timestamp 1666464484
transform 1 0 69104 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_669
timestamp 1666464484
transform 1 0 76272 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_673
timestamp 1666464484
transform 1 0 76720 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_676
timestamp 1666464484
transform 1 0 77056 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_740
timestamp 1666464484
transform 1 0 84224 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_744
timestamp 1666464484
transform 1 0 84672 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_747
timestamp 1666464484
transform 1 0 85008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_811
timestamp 1666464484
transform 1 0 92176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_815
timestamp 1666464484
transform 1 0 92624 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_818
timestamp 1666464484
transform 1 0 92960 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_882
timestamp 1666464484
transform 1 0 100128 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_886
timestamp 1666464484
transform 1 0 100576 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_889
timestamp 1666464484
transform 1 0 100912 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_953
timestamp 1666464484
transform 1 0 108080 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_957
timestamp 1666464484
transform 1 0 108528 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_960
timestamp 1666464484
transform 1 0 108864 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1024
timestamp 1666464484
transform 1 0 116032 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1028
timestamp 1666464484
transform 1 0 116480 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_1031
timestamp 1666464484
transform 1 0 116816 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1095
timestamp 1666464484
transform 1 0 123984 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1099
timestamp 1666464484
transform 1 0 124432 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_1102
timestamp 1666464484
transform 1 0 124768 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1166
timestamp 1666464484
transform 1 0 131936 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1170
timestamp 1666464484
transform 1 0 132384 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_1173
timestamp 1666464484
transform 1 0 132720 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1237
timestamp 1666464484
transform 1 0 139888 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1241
timestamp 1666464484
transform 1 0 140336 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_1244
timestamp 1666464484
transform 1 0 140672 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1308
timestamp 1666464484
transform 1 0 147840 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1312
timestamp 1666464484
transform 1 0 148288 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_1315
timestamp 1666464484
transform 1 0 148624 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1379
timestamp 1666464484
transform 1 0 155792 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1383
timestamp 1666464484
transform 1 0 156240 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_1386
timestamp 1666464484
transform 1 0 156576 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1450
timestamp 1666464484
transform 1 0 163744 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1454
timestamp 1666464484
transform 1 0 164192 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_1457
timestamp 1666464484
transform 1 0 164528 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1521
timestamp 1666464484
transform 1 0 171696 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1525
timestamp 1666464484
transform 1 0 172144 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_1528
timestamp 1666464484
transform 1 0 172480 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_90_1560
timestamp 1666464484
transform 1 0 176064 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1576
timestamp 1666464484
transform 1 0 177856 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1580
timestamp 1666464484
transform 1 0 178304 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_2
timestamp 1666464484
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_66
timestamp 1666464484
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_70
timestamp 1666464484
transform 1 0 9184 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_73
timestamp 1666464484
transform 1 0 9520 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_137
timestamp 1666464484
transform 1 0 16688 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_141
timestamp 1666464484
transform 1 0 17136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_144
timestamp 1666464484
transform 1 0 17472 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_208
timestamp 1666464484
transform 1 0 24640 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_212
timestamp 1666464484
transform 1 0 25088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_215
timestamp 1666464484
transform 1 0 25424 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_279
timestamp 1666464484
transform 1 0 32592 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_283
timestamp 1666464484
transform 1 0 33040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_286
timestamp 1666464484
transform 1 0 33376 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_350
timestamp 1666464484
transform 1 0 40544 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_354
timestamp 1666464484
transform 1 0 40992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_357
timestamp 1666464484
transform 1 0 41328 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_421
timestamp 1666464484
transform 1 0 48496 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_425
timestamp 1666464484
transform 1 0 48944 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_428
timestamp 1666464484
transform 1 0 49280 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_492
timestamp 1666464484
transform 1 0 56448 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_496
timestamp 1666464484
transform 1 0 56896 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_499
timestamp 1666464484
transform 1 0 57232 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_563
timestamp 1666464484
transform 1 0 64400 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_567
timestamp 1666464484
transform 1 0 64848 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_570
timestamp 1666464484
transform 1 0 65184 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_634
timestamp 1666464484
transform 1 0 72352 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_638
timestamp 1666464484
transform 1 0 72800 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_641
timestamp 1666464484
transform 1 0 73136 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_705
timestamp 1666464484
transform 1 0 80304 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_709
timestamp 1666464484
transform 1 0 80752 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_712
timestamp 1666464484
transform 1 0 81088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_776
timestamp 1666464484
transform 1 0 88256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_780
timestamp 1666464484
transform 1 0 88704 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_783
timestamp 1666464484
transform 1 0 89040 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_847
timestamp 1666464484
transform 1 0 96208 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_851
timestamp 1666464484
transform 1 0 96656 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_854
timestamp 1666464484
transform 1 0 96992 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_918
timestamp 1666464484
transform 1 0 104160 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_922
timestamp 1666464484
transform 1 0 104608 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_925
timestamp 1666464484
transform 1 0 104944 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_989
timestamp 1666464484
transform 1 0 112112 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_993
timestamp 1666464484
transform 1 0 112560 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_996
timestamp 1666464484
transform 1 0 112896 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_1060
timestamp 1666464484
transform 1 0 120064 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1064
timestamp 1666464484
transform 1 0 120512 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_1067
timestamp 1666464484
transform 1 0 120848 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_1131
timestamp 1666464484
transform 1 0 128016 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1135
timestamp 1666464484
transform 1 0 128464 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_1138
timestamp 1666464484
transform 1 0 128800 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_1202
timestamp 1666464484
transform 1 0 135968 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1206
timestamp 1666464484
transform 1 0 136416 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_1209
timestamp 1666464484
transform 1 0 136752 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_1273
timestamp 1666464484
transform 1 0 143920 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1277
timestamp 1666464484
transform 1 0 144368 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_1280
timestamp 1666464484
transform 1 0 144704 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_1344
timestamp 1666464484
transform 1 0 151872 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1348
timestamp 1666464484
transform 1 0 152320 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_1351
timestamp 1666464484
transform 1 0 152656 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_1415
timestamp 1666464484
transform 1 0 159824 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1419
timestamp 1666464484
transform 1 0 160272 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_1422
timestamp 1666464484
transform 1 0 160608 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_1486
timestamp 1666464484
transform 1 0 167776 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1490
timestamp 1666464484
transform 1 0 168224 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_1493
timestamp 1666464484
transform 1 0 168560 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_1557
timestamp 1666464484
transform 1 0 175728 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1561
timestamp 1666464484
transform 1 0 176176 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_1564
timestamp 1666464484
transform 1 0 176512 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1580
timestamp 1666464484
transform 1 0 178304 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_2
timestamp 1666464484
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_34
timestamp 1666464484
transform 1 0 5152 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_37
timestamp 1666464484
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_101
timestamp 1666464484
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_105
timestamp 1666464484
transform 1 0 13104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_108
timestamp 1666464484
transform 1 0 13440 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_172
timestamp 1666464484
transform 1 0 20608 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_176
timestamp 1666464484
transform 1 0 21056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_179
timestamp 1666464484
transform 1 0 21392 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_243
timestamp 1666464484
transform 1 0 28560 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_247
timestamp 1666464484
transform 1 0 29008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_250
timestamp 1666464484
transform 1 0 29344 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_314
timestamp 1666464484
transform 1 0 36512 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_318
timestamp 1666464484
transform 1 0 36960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_321
timestamp 1666464484
transform 1 0 37296 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_385
timestamp 1666464484
transform 1 0 44464 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_389
timestamp 1666464484
transform 1 0 44912 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_392
timestamp 1666464484
transform 1 0 45248 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_456
timestamp 1666464484
transform 1 0 52416 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_460
timestamp 1666464484
transform 1 0 52864 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_463
timestamp 1666464484
transform 1 0 53200 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_527
timestamp 1666464484
transform 1 0 60368 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_531
timestamp 1666464484
transform 1 0 60816 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_534
timestamp 1666464484
transform 1 0 61152 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_598
timestamp 1666464484
transform 1 0 68320 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_602
timestamp 1666464484
transform 1 0 68768 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_605
timestamp 1666464484
transform 1 0 69104 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_669
timestamp 1666464484
transform 1 0 76272 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_673
timestamp 1666464484
transform 1 0 76720 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_676
timestamp 1666464484
transform 1 0 77056 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_740
timestamp 1666464484
transform 1 0 84224 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_744
timestamp 1666464484
transform 1 0 84672 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_747
timestamp 1666464484
transform 1 0 85008 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_811
timestamp 1666464484
transform 1 0 92176 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_815
timestamp 1666464484
transform 1 0 92624 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_818
timestamp 1666464484
transform 1 0 92960 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_882
timestamp 1666464484
transform 1 0 100128 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_886
timestamp 1666464484
transform 1 0 100576 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_889
timestamp 1666464484
transform 1 0 100912 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_953
timestamp 1666464484
transform 1 0 108080 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_957
timestamp 1666464484
transform 1 0 108528 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_960
timestamp 1666464484
transform 1 0 108864 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1024
timestamp 1666464484
transform 1 0 116032 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1028
timestamp 1666464484
transform 1 0 116480 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_1031
timestamp 1666464484
transform 1 0 116816 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1095
timestamp 1666464484
transform 1 0 123984 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1099
timestamp 1666464484
transform 1 0 124432 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_1102
timestamp 1666464484
transform 1 0 124768 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1166
timestamp 1666464484
transform 1 0 131936 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1170
timestamp 1666464484
transform 1 0 132384 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_1173
timestamp 1666464484
transform 1 0 132720 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1237
timestamp 1666464484
transform 1 0 139888 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1241
timestamp 1666464484
transform 1 0 140336 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_1244
timestamp 1666464484
transform 1 0 140672 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1308
timestamp 1666464484
transform 1 0 147840 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1312
timestamp 1666464484
transform 1 0 148288 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_1315
timestamp 1666464484
transform 1 0 148624 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1379
timestamp 1666464484
transform 1 0 155792 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1383
timestamp 1666464484
transform 1 0 156240 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_1386
timestamp 1666464484
transform 1 0 156576 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1450
timestamp 1666464484
transform 1 0 163744 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1454
timestamp 1666464484
transform 1 0 164192 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_1457
timestamp 1666464484
transform 1 0 164528 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1521
timestamp 1666464484
transform 1 0 171696 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1525
timestamp 1666464484
transform 1 0 172144 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_1528
timestamp 1666464484
transform 1 0 172480 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_1560
timestamp 1666464484
transform 1 0 176064 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1576
timestamp 1666464484
transform 1 0 177856 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1580
timestamp 1666464484
transform 1 0 178304 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_2
timestamp 1666464484
transform 1 0 1568 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_66
timestamp 1666464484
transform 1 0 8736 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_70
timestamp 1666464484
transform 1 0 9184 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_73
timestamp 1666464484
transform 1 0 9520 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_137
timestamp 1666464484
transform 1 0 16688 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_141
timestamp 1666464484
transform 1 0 17136 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_144
timestamp 1666464484
transform 1 0 17472 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_208
timestamp 1666464484
transform 1 0 24640 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_212
timestamp 1666464484
transform 1 0 25088 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_215
timestamp 1666464484
transform 1 0 25424 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_279
timestamp 1666464484
transform 1 0 32592 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_283
timestamp 1666464484
transform 1 0 33040 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_286
timestamp 1666464484
transform 1 0 33376 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_350
timestamp 1666464484
transform 1 0 40544 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_354
timestamp 1666464484
transform 1 0 40992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_357
timestamp 1666464484
transform 1 0 41328 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_421
timestamp 1666464484
transform 1 0 48496 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_425
timestamp 1666464484
transform 1 0 48944 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_428
timestamp 1666464484
transform 1 0 49280 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_492
timestamp 1666464484
transform 1 0 56448 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_496
timestamp 1666464484
transform 1 0 56896 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_499
timestamp 1666464484
transform 1 0 57232 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_563
timestamp 1666464484
transform 1 0 64400 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_567
timestamp 1666464484
transform 1 0 64848 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_570
timestamp 1666464484
transform 1 0 65184 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_634
timestamp 1666464484
transform 1 0 72352 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_638
timestamp 1666464484
transform 1 0 72800 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_641
timestamp 1666464484
transform 1 0 73136 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_705
timestamp 1666464484
transform 1 0 80304 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_709
timestamp 1666464484
transform 1 0 80752 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_712
timestamp 1666464484
transform 1 0 81088 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_776
timestamp 1666464484
transform 1 0 88256 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_780
timestamp 1666464484
transform 1 0 88704 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_783
timestamp 1666464484
transform 1 0 89040 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_847
timestamp 1666464484
transform 1 0 96208 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_851
timestamp 1666464484
transform 1 0 96656 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_854
timestamp 1666464484
transform 1 0 96992 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_918
timestamp 1666464484
transform 1 0 104160 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_922
timestamp 1666464484
transform 1 0 104608 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_925
timestamp 1666464484
transform 1 0 104944 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_989
timestamp 1666464484
transform 1 0 112112 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_993
timestamp 1666464484
transform 1 0 112560 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_996
timestamp 1666464484
transform 1 0 112896 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_1060
timestamp 1666464484
transform 1 0 120064 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1064
timestamp 1666464484
transform 1 0 120512 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_1067
timestamp 1666464484
transform 1 0 120848 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_1131
timestamp 1666464484
transform 1 0 128016 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1135
timestamp 1666464484
transform 1 0 128464 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_1138
timestamp 1666464484
transform 1 0 128800 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_1202
timestamp 1666464484
transform 1 0 135968 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1206
timestamp 1666464484
transform 1 0 136416 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_1209
timestamp 1666464484
transform 1 0 136752 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_1273
timestamp 1666464484
transform 1 0 143920 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1277
timestamp 1666464484
transform 1 0 144368 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_1280
timestamp 1666464484
transform 1 0 144704 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_1344
timestamp 1666464484
transform 1 0 151872 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1348
timestamp 1666464484
transform 1 0 152320 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_1351
timestamp 1666464484
transform 1 0 152656 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_1415
timestamp 1666464484
transform 1 0 159824 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1419
timestamp 1666464484
transform 1 0 160272 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_1422
timestamp 1666464484
transform 1 0 160608 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_1486
timestamp 1666464484
transform 1 0 167776 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1490
timestamp 1666464484
transform 1 0 168224 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_1493
timestamp 1666464484
transform 1 0 168560 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_1557
timestamp 1666464484
transform 1 0 175728 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1561
timestamp 1666464484
transform 1 0 176176 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_1564
timestamp 1666464484
transform 1 0 176512 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1580
timestamp 1666464484
transform 1 0 178304 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_94_2
timestamp 1666464484
transform 1 0 1568 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_34
timestamp 1666464484
transform 1 0 5152 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_37
timestamp 1666464484
transform 1 0 5488 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_101
timestamp 1666464484
transform 1 0 12656 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_105
timestamp 1666464484
transform 1 0 13104 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_108
timestamp 1666464484
transform 1 0 13440 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_172
timestamp 1666464484
transform 1 0 20608 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_176
timestamp 1666464484
transform 1 0 21056 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_179
timestamp 1666464484
transform 1 0 21392 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_243
timestamp 1666464484
transform 1 0 28560 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_247
timestamp 1666464484
transform 1 0 29008 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_250
timestamp 1666464484
transform 1 0 29344 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_314
timestamp 1666464484
transform 1 0 36512 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_318
timestamp 1666464484
transform 1 0 36960 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_321
timestamp 1666464484
transform 1 0 37296 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_385
timestamp 1666464484
transform 1 0 44464 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_389
timestamp 1666464484
transform 1 0 44912 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_392
timestamp 1666464484
transform 1 0 45248 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_456
timestamp 1666464484
transform 1 0 52416 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_460
timestamp 1666464484
transform 1 0 52864 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_463
timestamp 1666464484
transform 1 0 53200 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_527
timestamp 1666464484
transform 1 0 60368 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_531
timestamp 1666464484
transform 1 0 60816 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_534
timestamp 1666464484
transform 1 0 61152 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_598
timestamp 1666464484
transform 1 0 68320 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_602
timestamp 1666464484
transform 1 0 68768 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_605
timestamp 1666464484
transform 1 0 69104 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_669
timestamp 1666464484
transform 1 0 76272 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_673
timestamp 1666464484
transform 1 0 76720 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_676
timestamp 1666464484
transform 1 0 77056 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_740
timestamp 1666464484
transform 1 0 84224 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_744
timestamp 1666464484
transform 1 0 84672 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_747
timestamp 1666464484
transform 1 0 85008 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_811
timestamp 1666464484
transform 1 0 92176 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_815
timestamp 1666464484
transform 1 0 92624 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_818
timestamp 1666464484
transform 1 0 92960 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_882
timestamp 1666464484
transform 1 0 100128 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_886
timestamp 1666464484
transform 1 0 100576 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_889
timestamp 1666464484
transform 1 0 100912 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_953
timestamp 1666464484
transform 1 0 108080 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_957
timestamp 1666464484
transform 1 0 108528 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_960
timestamp 1666464484
transform 1 0 108864 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1024
timestamp 1666464484
transform 1 0 116032 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1028
timestamp 1666464484
transform 1 0 116480 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_1031
timestamp 1666464484
transform 1 0 116816 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1095
timestamp 1666464484
transform 1 0 123984 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1099
timestamp 1666464484
transform 1 0 124432 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_1102
timestamp 1666464484
transform 1 0 124768 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1166
timestamp 1666464484
transform 1 0 131936 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1170
timestamp 1666464484
transform 1 0 132384 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_1173
timestamp 1666464484
transform 1 0 132720 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1237
timestamp 1666464484
transform 1 0 139888 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1241
timestamp 1666464484
transform 1 0 140336 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_1244
timestamp 1666464484
transform 1 0 140672 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1308
timestamp 1666464484
transform 1 0 147840 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1312
timestamp 1666464484
transform 1 0 148288 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_1315
timestamp 1666464484
transform 1 0 148624 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1379
timestamp 1666464484
transform 1 0 155792 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1383
timestamp 1666464484
transform 1 0 156240 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_1386
timestamp 1666464484
transform 1 0 156576 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1450
timestamp 1666464484
transform 1 0 163744 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1454
timestamp 1666464484
transform 1 0 164192 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_1457
timestamp 1666464484
transform 1 0 164528 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1521
timestamp 1666464484
transform 1 0 171696 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1525
timestamp 1666464484
transform 1 0 172144 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_94_1528
timestamp 1666464484
transform 1 0 172480 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_94_1560
timestamp 1666464484
transform 1 0 176064 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1576
timestamp 1666464484
transform 1 0 177856 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1580
timestamp 1666464484
transform 1 0 178304 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_2
timestamp 1666464484
transform 1 0 1568 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_66
timestamp 1666464484
transform 1 0 8736 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_70
timestamp 1666464484
transform 1 0 9184 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_73
timestamp 1666464484
transform 1 0 9520 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_137
timestamp 1666464484
transform 1 0 16688 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_141
timestamp 1666464484
transform 1 0 17136 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_144
timestamp 1666464484
transform 1 0 17472 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_208
timestamp 1666464484
transform 1 0 24640 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_212
timestamp 1666464484
transform 1 0 25088 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_215
timestamp 1666464484
transform 1 0 25424 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_279
timestamp 1666464484
transform 1 0 32592 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_283
timestamp 1666464484
transform 1 0 33040 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_286
timestamp 1666464484
transform 1 0 33376 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_350
timestamp 1666464484
transform 1 0 40544 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_354
timestamp 1666464484
transform 1 0 40992 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_357
timestamp 1666464484
transform 1 0 41328 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_421
timestamp 1666464484
transform 1 0 48496 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_425
timestamp 1666464484
transform 1 0 48944 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_428
timestamp 1666464484
transform 1 0 49280 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_492
timestamp 1666464484
transform 1 0 56448 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_496
timestamp 1666464484
transform 1 0 56896 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_499
timestamp 1666464484
transform 1 0 57232 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_563
timestamp 1666464484
transform 1 0 64400 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_567
timestamp 1666464484
transform 1 0 64848 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_570
timestamp 1666464484
transform 1 0 65184 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_634
timestamp 1666464484
transform 1 0 72352 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_638
timestamp 1666464484
transform 1 0 72800 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_641
timestamp 1666464484
transform 1 0 73136 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_705
timestamp 1666464484
transform 1 0 80304 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_709
timestamp 1666464484
transform 1 0 80752 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_712
timestamp 1666464484
transform 1 0 81088 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_776
timestamp 1666464484
transform 1 0 88256 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_780
timestamp 1666464484
transform 1 0 88704 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_783
timestamp 1666464484
transform 1 0 89040 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_847
timestamp 1666464484
transform 1 0 96208 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_851
timestamp 1666464484
transform 1 0 96656 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_854
timestamp 1666464484
transform 1 0 96992 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_918
timestamp 1666464484
transform 1 0 104160 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_922
timestamp 1666464484
transform 1 0 104608 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_925
timestamp 1666464484
transform 1 0 104944 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_989
timestamp 1666464484
transform 1 0 112112 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_993
timestamp 1666464484
transform 1 0 112560 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_996
timestamp 1666464484
transform 1 0 112896 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_1060
timestamp 1666464484
transform 1 0 120064 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1064
timestamp 1666464484
transform 1 0 120512 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_1067
timestamp 1666464484
transform 1 0 120848 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_1131
timestamp 1666464484
transform 1 0 128016 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1135
timestamp 1666464484
transform 1 0 128464 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_1138
timestamp 1666464484
transform 1 0 128800 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_1202
timestamp 1666464484
transform 1 0 135968 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1206
timestamp 1666464484
transform 1 0 136416 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_1209
timestamp 1666464484
transform 1 0 136752 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_1273
timestamp 1666464484
transform 1 0 143920 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1277
timestamp 1666464484
transform 1 0 144368 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_1280
timestamp 1666464484
transform 1 0 144704 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_1344
timestamp 1666464484
transform 1 0 151872 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1348
timestamp 1666464484
transform 1 0 152320 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_1351
timestamp 1666464484
transform 1 0 152656 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_1415
timestamp 1666464484
transform 1 0 159824 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1419
timestamp 1666464484
transform 1 0 160272 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_1422
timestamp 1666464484
transform 1 0 160608 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_1486
timestamp 1666464484
transform 1 0 167776 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1490
timestamp 1666464484
transform 1 0 168224 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_1493
timestamp 1666464484
transform 1 0 168560 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_1557
timestamp 1666464484
transform 1 0 175728 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1561
timestamp 1666464484
transform 1 0 176176 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_95_1564
timestamp 1666464484
transform 1 0 176512 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1580
timestamp 1666464484
transform 1 0 178304 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_96_2
timestamp 1666464484
transform 1 0 1568 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_34
timestamp 1666464484
transform 1 0 5152 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_37
timestamp 1666464484
transform 1 0 5488 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_101
timestamp 1666464484
transform 1 0 12656 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_105
timestamp 1666464484
transform 1 0 13104 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_108
timestamp 1666464484
transform 1 0 13440 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_172
timestamp 1666464484
transform 1 0 20608 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_176
timestamp 1666464484
transform 1 0 21056 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_179
timestamp 1666464484
transform 1 0 21392 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_243
timestamp 1666464484
transform 1 0 28560 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_247
timestamp 1666464484
transform 1 0 29008 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_250
timestamp 1666464484
transform 1 0 29344 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_314
timestamp 1666464484
transform 1 0 36512 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_318
timestamp 1666464484
transform 1 0 36960 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_321
timestamp 1666464484
transform 1 0 37296 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_385
timestamp 1666464484
transform 1 0 44464 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_389
timestamp 1666464484
transform 1 0 44912 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_392
timestamp 1666464484
transform 1 0 45248 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_456
timestamp 1666464484
transform 1 0 52416 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_460
timestamp 1666464484
transform 1 0 52864 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_463
timestamp 1666464484
transform 1 0 53200 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_527
timestamp 1666464484
transform 1 0 60368 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_531
timestamp 1666464484
transform 1 0 60816 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_534
timestamp 1666464484
transform 1 0 61152 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_598
timestamp 1666464484
transform 1 0 68320 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_602
timestamp 1666464484
transform 1 0 68768 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_605
timestamp 1666464484
transform 1 0 69104 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_669
timestamp 1666464484
transform 1 0 76272 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_673
timestamp 1666464484
transform 1 0 76720 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_676
timestamp 1666464484
transform 1 0 77056 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_740
timestamp 1666464484
transform 1 0 84224 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_744
timestamp 1666464484
transform 1 0 84672 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_747
timestamp 1666464484
transform 1 0 85008 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_811
timestamp 1666464484
transform 1 0 92176 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_815
timestamp 1666464484
transform 1 0 92624 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_818
timestamp 1666464484
transform 1 0 92960 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_882
timestamp 1666464484
transform 1 0 100128 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_886
timestamp 1666464484
transform 1 0 100576 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_889
timestamp 1666464484
transform 1 0 100912 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_953
timestamp 1666464484
transform 1 0 108080 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_957
timestamp 1666464484
transform 1 0 108528 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_960
timestamp 1666464484
transform 1 0 108864 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1024
timestamp 1666464484
transform 1 0 116032 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1028
timestamp 1666464484
transform 1 0 116480 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_1031
timestamp 1666464484
transform 1 0 116816 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1095
timestamp 1666464484
transform 1 0 123984 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1099
timestamp 1666464484
transform 1 0 124432 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_1102
timestamp 1666464484
transform 1 0 124768 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1166
timestamp 1666464484
transform 1 0 131936 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1170
timestamp 1666464484
transform 1 0 132384 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_1173
timestamp 1666464484
transform 1 0 132720 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1237
timestamp 1666464484
transform 1 0 139888 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1241
timestamp 1666464484
transform 1 0 140336 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_1244
timestamp 1666464484
transform 1 0 140672 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1308
timestamp 1666464484
transform 1 0 147840 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1312
timestamp 1666464484
transform 1 0 148288 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_1315
timestamp 1666464484
transform 1 0 148624 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1379
timestamp 1666464484
transform 1 0 155792 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1383
timestamp 1666464484
transform 1 0 156240 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_1386
timestamp 1666464484
transform 1 0 156576 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1450
timestamp 1666464484
transform 1 0 163744 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1454
timestamp 1666464484
transform 1 0 164192 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_1457
timestamp 1666464484
transform 1 0 164528 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1521
timestamp 1666464484
transform 1 0 171696 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1525
timestamp 1666464484
transform 1 0 172144 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_96_1528
timestamp 1666464484
transform 1 0 172480 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_96_1560
timestamp 1666464484
transform 1 0 176064 0 1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1576
timestamp 1666464484
transform 1 0 177856 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1580
timestamp 1666464484
transform 1 0 178304 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_2
timestamp 1666464484
transform 1 0 1568 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_66
timestamp 1666464484
transform 1 0 8736 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_70
timestamp 1666464484
transform 1 0 9184 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_73
timestamp 1666464484
transform 1 0 9520 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_137
timestamp 1666464484
transform 1 0 16688 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_141
timestamp 1666464484
transform 1 0 17136 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_144
timestamp 1666464484
transform 1 0 17472 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_208
timestamp 1666464484
transform 1 0 24640 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_212
timestamp 1666464484
transform 1 0 25088 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_215
timestamp 1666464484
transform 1 0 25424 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_279
timestamp 1666464484
transform 1 0 32592 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_283
timestamp 1666464484
transform 1 0 33040 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_286
timestamp 1666464484
transform 1 0 33376 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_350
timestamp 1666464484
transform 1 0 40544 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_354
timestamp 1666464484
transform 1 0 40992 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_357
timestamp 1666464484
transform 1 0 41328 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_421
timestamp 1666464484
transform 1 0 48496 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_425
timestamp 1666464484
transform 1 0 48944 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_428
timestamp 1666464484
transform 1 0 49280 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_492
timestamp 1666464484
transform 1 0 56448 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_496
timestamp 1666464484
transform 1 0 56896 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_499
timestamp 1666464484
transform 1 0 57232 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_563
timestamp 1666464484
transform 1 0 64400 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_567
timestamp 1666464484
transform 1 0 64848 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_570
timestamp 1666464484
transform 1 0 65184 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_634
timestamp 1666464484
transform 1 0 72352 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_638
timestamp 1666464484
transform 1 0 72800 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_641
timestamp 1666464484
transform 1 0 73136 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_705
timestamp 1666464484
transform 1 0 80304 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_709
timestamp 1666464484
transform 1 0 80752 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_712
timestamp 1666464484
transform 1 0 81088 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_776
timestamp 1666464484
transform 1 0 88256 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_780
timestamp 1666464484
transform 1 0 88704 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_783
timestamp 1666464484
transform 1 0 89040 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_847
timestamp 1666464484
transform 1 0 96208 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_851
timestamp 1666464484
transform 1 0 96656 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_854
timestamp 1666464484
transform 1 0 96992 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_918
timestamp 1666464484
transform 1 0 104160 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_922
timestamp 1666464484
transform 1 0 104608 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_925
timestamp 1666464484
transform 1 0 104944 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_989
timestamp 1666464484
transform 1 0 112112 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_993
timestamp 1666464484
transform 1 0 112560 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_996
timestamp 1666464484
transform 1 0 112896 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1060
timestamp 1666464484
transform 1 0 120064 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1064
timestamp 1666464484
transform 1 0 120512 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_1067
timestamp 1666464484
transform 1 0 120848 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1131
timestamp 1666464484
transform 1 0 128016 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1135
timestamp 1666464484
transform 1 0 128464 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_1138
timestamp 1666464484
transform 1 0 128800 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1202
timestamp 1666464484
transform 1 0 135968 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1206
timestamp 1666464484
transform 1 0 136416 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_1209
timestamp 1666464484
transform 1 0 136752 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1273
timestamp 1666464484
transform 1 0 143920 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1277
timestamp 1666464484
transform 1 0 144368 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_1280
timestamp 1666464484
transform 1 0 144704 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1344
timestamp 1666464484
transform 1 0 151872 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1348
timestamp 1666464484
transform 1 0 152320 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_1351
timestamp 1666464484
transform 1 0 152656 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1415
timestamp 1666464484
transform 1 0 159824 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1419
timestamp 1666464484
transform 1 0 160272 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_1422
timestamp 1666464484
transform 1 0 160608 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1486
timestamp 1666464484
transform 1 0 167776 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1490
timestamp 1666464484
transform 1 0 168224 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_1493
timestamp 1666464484
transform 1 0 168560 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1557
timestamp 1666464484
transform 1 0 175728 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1561
timestamp 1666464484
transform 1 0 176176 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_97_1564
timestamp 1666464484
transform 1 0 176512 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1580
timestamp 1666464484
transform 1 0 178304 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_98_2
timestamp 1666464484
transform 1 0 1568 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_34
timestamp 1666464484
transform 1 0 5152 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_37
timestamp 1666464484
transform 1 0 5488 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_101
timestamp 1666464484
transform 1 0 12656 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_105
timestamp 1666464484
transform 1 0 13104 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_108
timestamp 1666464484
transform 1 0 13440 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_172
timestamp 1666464484
transform 1 0 20608 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_176
timestamp 1666464484
transform 1 0 21056 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_179
timestamp 1666464484
transform 1 0 21392 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_243
timestamp 1666464484
transform 1 0 28560 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_247
timestamp 1666464484
transform 1 0 29008 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_250
timestamp 1666464484
transform 1 0 29344 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_314
timestamp 1666464484
transform 1 0 36512 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_318
timestamp 1666464484
transform 1 0 36960 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_321
timestamp 1666464484
transform 1 0 37296 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_385
timestamp 1666464484
transform 1 0 44464 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_389
timestamp 1666464484
transform 1 0 44912 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_392
timestamp 1666464484
transform 1 0 45248 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_456
timestamp 1666464484
transform 1 0 52416 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_460
timestamp 1666464484
transform 1 0 52864 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_463
timestamp 1666464484
transform 1 0 53200 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_527
timestamp 1666464484
transform 1 0 60368 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_531
timestamp 1666464484
transform 1 0 60816 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_534
timestamp 1666464484
transform 1 0 61152 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_598
timestamp 1666464484
transform 1 0 68320 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_602
timestamp 1666464484
transform 1 0 68768 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_605
timestamp 1666464484
transform 1 0 69104 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_669
timestamp 1666464484
transform 1 0 76272 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_673
timestamp 1666464484
transform 1 0 76720 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_676
timestamp 1666464484
transform 1 0 77056 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_740
timestamp 1666464484
transform 1 0 84224 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_744
timestamp 1666464484
transform 1 0 84672 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_747
timestamp 1666464484
transform 1 0 85008 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_811
timestamp 1666464484
transform 1 0 92176 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_815
timestamp 1666464484
transform 1 0 92624 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_818
timestamp 1666464484
transform 1 0 92960 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_882
timestamp 1666464484
transform 1 0 100128 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_886
timestamp 1666464484
transform 1 0 100576 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_889
timestamp 1666464484
transform 1 0 100912 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_953
timestamp 1666464484
transform 1 0 108080 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_957
timestamp 1666464484
transform 1 0 108528 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_960
timestamp 1666464484
transform 1 0 108864 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1024
timestamp 1666464484
transform 1 0 116032 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1028
timestamp 1666464484
transform 1 0 116480 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_1031
timestamp 1666464484
transform 1 0 116816 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1095
timestamp 1666464484
transform 1 0 123984 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1099
timestamp 1666464484
transform 1 0 124432 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_1102
timestamp 1666464484
transform 1 0 124768 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1166
timestamp 1666464484
transform 1 0 131936 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1170
timestamp 1666464484
transform 1 0 132384 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_1173
timestamp 1666464484
transform 1 0 132720 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1237
timestamp 1666464484
transform 1 0 139888 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1241
timestamp 1666464484
transform 1 0 140336 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_1244
timestamp 1666464484
transform 1 0 140672 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1308
timestamp 1666464484
transform 1 0 147840 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1312
timestamp 1666464484
transform 1 0 148288 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_1315
timestamp 1666464484
transform 1 0 148624 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1379
timestamp 1666464484
transform 1 0 155792 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1383
timestamp 1666464484
transform 1 0 156240 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_1386
timestamp 1666464484
transform 1 0 156576 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1450
timestamp 1666464484
transform 1 0 163744 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1454
timestamp 1666464484
transform 1 0 164192 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_1457
timestamp 1666464484
transform 1 0 164528 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1521
timestamp 1666464484
transform 1 0 171696 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1525
timestamp 1666464484
transform 1 0 172144 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_98_1528
timestamp 1666464484
transform 1 0 172480 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_98_1560
timestamp 1666464484
transform 1 0 176064 0 1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1576
timestamp 1666464484
transform 1 0 177856 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1580
timestamp 1666464484
transform 1 0 178304 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_2
timestamp 1666464484
transform 1 0 1568 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_66
timestamp 1666464484
transform 1 0 8736 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_70
timestamp 1666464484
transform 1 0 9184 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_73
timestamp 1666464484
transform 1 0 9520 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_137
timestamp 1666464484
transform 1 0 16688 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_141
timestamp 1666464484
transform 1 0 17136 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_144
timestamp 1666464484
transform 1 0 17472 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_208
timestamp 1666464484
transform 1 0 24640 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_212
timestamp 1666464484
transform 1 0 25088 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_215
timestamp 1666464484
transform 1 0 25424 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_279
timestamp 1666464484
transform 1 0 32592 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_283
timestamp 1666464484
transform 1 0 33040 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_286
timestamp 1666464484
transform 1 0 33376 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_350
timestamp 1666464484
transform 1 0 40544 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_354
timestamp 1666464484
transform 1 0 40992 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_357
timestamp 1666464484
transform 1 0 41328 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_421
timestamp 1666464484
transform 1 0 48496 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_425
timestamp 1666464484
transform 1 0 48944 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_428
timestamp 1666464484
transform 1 0 49280 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_492
timestamp 1666464484
transform 1 0 56448 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_496
timestamp 1666464484
transform 1 0 56896 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_499
timestamp 1666464484
transform 1 0 57232 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_563
timestamp 1666464484
transform 1 0 64400 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_567
timestamp 1666464484
transform 1 0 64848 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_570
timestamp 1666464484
transform 1 0 65184 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_634
timestamp 1666464484
transform 1 0 72352 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_638
timestamp 1666464484
transform 1 0 72800 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_641
timestamp 1666464484
transform 1 0 73136 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_705
timestamp 1666464484
transform 1 0 80304 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_709
timestamp 1666464484
transform 1 0 80752 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_712
timestamp 1666464484
transform 1 0 81088 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_776
timestamp 1666464484
transform 1 0 88256 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_780
timestamp 1666464484
transform 1 0 88704 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_783
timestamp 1666464484
transform 1 0 89040 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_847
timestamp 1666464484
transform 1 0 96208 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_851
timestamp 1666464484
transform 1 0 96656 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_854
timestamp 1666464484
transform 1 0 96992 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_918
timestamp 1666464484
transform 1 0 104160 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_922
timestamp 1666464484
transform 1 0 104608 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_925
timestamp 1666464484
transform 1 0 104944 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_989
timestamp 1666464484
transform 1 0 112112 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_993
timestamp 1666464484
transform 1 0 112560 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_996
timestamp 1666464484
transform 1 0 112896 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_1060
timestamp 1666464484
transform 1 0 120064 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1064
timestamp 1666464484
transform 1 0 120512 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_1067
timestamp 1666464484
transform 1 0 120848 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_1131
timestamp 1666464484
transform 1 0 128016 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1135
timestamp 1666464484
transform 1 0 128464 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_1138
timestamp 1666464484
transform 1 0 128800 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_1202
timestamp 1666464484
transform 1 0 135968 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1206
timestamp 1666464484
transform 1 0 136416 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_1209
timestamp 1666464484
transform 1 0 136752 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_1273
timestamp 1666464484
transform 1 0 143920 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1277
timestamp 1666464484
transform 1 0 144368 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_1280
timestamp 1666464484
transform 1 0 144704 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_1344
timestamp 1666464484
transform 1 0 151872 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1348
timestamp 1666464484
transform 1 0 152320 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_1351
timestamp 1666464484
transform 1 0 152656 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_1415
timestamp 1666464484
transform 1 0 159824 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1419
timestamp 1666464484
transform 1 0 160272 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_1422
timestamp 1666464484
transform 1 0 160608 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_1486
timestamp 1666464484
transform 1 0 167776 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1490
timestamp 1666464484
transform 1 0 168224 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_1493
timestamp 1666464484
transform 1 0 168560 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_1557
timestamp 1666464484
transform 1 0 175728 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1561
timestamp 1666464484
transform 1 0 176176 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_99_1564
timestamp 1666464484
transform 1 0 176512 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1580
timestamp 1666464484
transform 1 0 178304 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_100_2
timestamp 1666464484
transform 1 0 1568 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_34
timestamp 1666464484
transform 1 0 5152 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_37
timestamp 1666464484
transform 1 0 5488 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_101
timestamp 1666464484
transform 1 0 12656 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_105
timestamp 1666464484
transform 1 0 13104 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_108
timestamp 1666464484
transform 1 0 13440 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_172
timestamp 1666464484
transform 1 0 20608 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_176
timestamp 1666464484
transform 1 0 21056 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_179
timestamp 1666464484
transform 1 0 21392 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_243
timestamp 1666464484
transform 1 0 28560 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_247
timestamp 1666464484
transform 1 0 29008 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_250
timestamp 1666464484
transform 1 0 29344 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_314
timestamp 1666464484
transform 1 0 36512 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_318
timestamp 1666464484
transform 1 0 36960 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_321
timestamp 1666464484
transform 1 0 37296 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_385
timestamp 1666464484
transform 1 0 44464 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_389
timestamp 1666464484
transform 1 0 44912 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_392
timestamp 1666464484
transform 1 0 45248 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_456
timestamp 1666464484
transform 1 0 52416 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_460
timestamp 1666464484
transform 1 0 52864 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_463
timestamp 1666464484
transform 1 0 53200 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_527
timestamp 1666464484
transform 1 0 60368 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_531
timestamp 1666464484
transform 1 0 60816 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_534
timestamp 1666464484
transform 1 0 61152 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_598
timestamp 1666464484
transform 1 0 68320 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_602
timestamp 1666464484
transform 1 0 68768 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_605
timestamp 1666464484
transform 1 0 69104 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_669
timestamp 1666464484
transform 1 0 76272 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_673
timestamp 1666464484
transform 1 0 76720 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_676
timestamp 1666464484
transform 1 0 77056 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_740
timestamp 1666464484
transform 1 0 84224 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_744
timestamp 1666464484
transform 1 0 84672 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_747
timestamp 1666464484
transform 1 0 85008 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_811
timestamp 1666464484
transform 1 0 92176 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_815
timestamp 1666464484
transform 1 0 92624 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_818
timestamp 1666464484
transform 1 0 92960 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_882
timestamp 1666464484
transform 1 0 100128 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_886
timestamp 1666464484
transform 1 0 100576 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_889
timestamp 1666464484
transform 1 0 100912 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_953
timestamp 1666464484
transform 1 0 108080 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_957
timestamp 1666464484
transform 1 0 108528 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_960
timestamp 1666464484
transform 1 0 108864 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1024
timestamp 1666464484
transform 1 0 116032 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1028
timestamp 1666464484
transform 1 0 116480 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_1031
timestamp 1666464484
transform 1 0 116816 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1095
timestamp 1666464484
transform 1 0 123984 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1099
timestamp 1666464484
transform 1 0 124432 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_1102
timestamp 1666464484
transform 1 0 124768 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1166
timestamp 1666464484
transform 1 0 131936 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1170
timestamp 1666464484
transform 1 0 132384 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_1173
timestamp 1666464484
transform 1 0 132720 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1237
timestamp 1666464484
transform 1 0 139888 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1241
timestamp 1666464484
transform 1 0 140336 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_1244
timestamp 1666464484
transform 1 0 140672 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1308
timestamp 1666464484
transform 1 0 147840 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1312
timestamp 1666464484
transform 1 0 148288 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_1315
timestamp 1666464484
transform 1 0 148624 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1379
timestamp 1666464484
transform 1 0 155792 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1383
timestamp 1666464484
transform 1 0 156240 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_1386
timestamp 1666464484
transform 1 0 156576 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1450
timestamp 1666464484
transform 1 0 163744 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1454
timestamp 1666464484
transform 1 0 164192 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_1457
timestamp 1666464484
transform 1 0 164528 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1521
timestamp 1666464484
transform 1 0 171696 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1525
timestamp 1666464484
transform 1 0 172144 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_100_1528
timestamp 1666464484
transform 1 0 172480 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_100_1560
timestamp 1666464484
transform 1 0 176064 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1576
timestamp 1666464484
transform 1 0 177856 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1580
timestamp 1666464484
transform 1 0 178304 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_2
timestamp 1666464484
transform 1 0 1568 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_66
timestamp 1666464484
transform 1 0 8736 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_70
timestamp 1666464484
transform 1 0 9184 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_73
timestamp 1666464484
transform 1 0 9520 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_137
timestamp 1666464484
transform 1 0 16688 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_141
timestamp 1666464484
transform 1 0 17136 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_144
timestamp 1666464484
transform 1 0 17472 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_208
timestamp 1666464484
transform 1 0 24640 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_212
timestamp 1666464484
transform 1 0 25088 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_215
timestamp 1666464484
transform 1 0 25424 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_279
timestamp 1666464484
transform 1 0 32592 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_283
timestamp 1666464484
transform 1 0 33040 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_286
timestamp 1666464484
transform 1 0 33376 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_350
timestamp 1666464484
transform 1 0 40544 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_354
timestamp 1666464484
transform 1 0 40992 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_357
timestamp 1666464484
transform 1 0 41328 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_421
timestamp 1666464484
transform 1 0 48496 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_425
timestamp 1666464484
transform 1 0 48944 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_428
timestamp 1666464484
transform 1 0 49280 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_492
timestamp 1666464484
transform 1 0 56448 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_496
timestamp 1666464484
transform 1 0 56896 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_499
timestamp 1666464484
transform 1 0 57232 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_563
timestamp 1666464484
transform 1 0 64400 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_567
timestamp 1666464484
transform 1 0 64848 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_570
timestamp 1666464484
transform 1 0 65184 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_634
timestamp 1666464484
transform 1 0 72352 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_638
timestamp 1666464484
transform 1 0 72800 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_641
timestamp 1666464484
transform 1 0 73136 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_705
timestamp 1666464484
transform 1 0 80304 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_709
timestamp 1666464484
transform 1 0 80752 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_712
timestamp 1666464484
transform 1 0 81088 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_776
timestamp 1666464484
transform 1 0 88256 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_780
timestamp 1666464484
transform 1 0 88704 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_783
timestamp 1666464484
transform 1 0 89040 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_847
timestamp 1666464484
transform 1 0 96208 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_851
timestamp 1666464484
transform 1 0 96656 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_854
timestamp 1666464484
transform 1 0 96992 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_918
timestamp 1666464484
transform 1 0 104160 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_922
timestamp 1666464484
transform 1 0 104608 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_925
timestamp 1666464484
transform 1 0 104944 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_989
timestamp 1666464484
transform 1 0 112112 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_993
timestamp 1666464484
transform 1 0 112560 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_996
timestamp 1666464484
transform 1 0 112896 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1060
timestamp 1666464484
transform 1 0 120064 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1064
timestamp 1666464484
transform 1 0 120512 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_1067
timestamp 1666464484
transform 1 0 120848 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1131
timestamp 1666464484
transform 1 0 128016 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1135
timestamp 1666464484
transform 1 0 128464 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_1138
timestamp 1666464484
transform 1 0 128800 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1202
timestamp 1666464484
transform 1 0 135968 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1206
timestamp 1666464484
transform 1 0 136416 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_1209
timestamp 1666464484
transform 1 0 136752 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1273
timestamp 1666464484
transform 1 0 143920 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1277
timestamp 1666464484
transform 1 0 144368 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_1280
timestamp 1666464484
transform 1 0 144704 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1344
timestamp 1666464484
transform 1 0 151872 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1348
timestamp 1666464484
transform 1 0 152320 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_1351
timestamp 1666464484
transform 1 0 152656 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1415
timestamp 1666464484
transform 1 0 159824 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1419
timestamp 1666464484
transform 1 0 160272 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_1422
timestamp 1666464484
transform 1 0 160608 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1486
timestamp 1666464484
transform 1 0 167776 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1490
timestamp 1666464484
transform 1 0 168224 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_1493
timestamp 1666464484
transform 1 0 168560 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1557
timestamp 1666464484
transform 1 0 175728 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1561
timestamp 1666464484
transform 1 0 176176 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_101_1564
timestamp 1666464484
transform 1 0 176512 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1580
timestamp 1666464484
transform 1 0 178304 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_102_2
timestamp 1666464484
transform 1 0 1568 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_34
timestamp 1666464484
transform 1 0 5152 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_37
timestamp 1666464484
transform 1 0 5488 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_101
timestamp 1666464484
transform 1 0 12656 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_105
timestamp 1666464484
transform 1 0 13104 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_108
timestamp 1666464484
transform 1 0 13440 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_172
timestamp 1666464484
transform 1 0 20608 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_176
timestamp 1666464484
transform 1 0 21056 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_179
timestamp 1666464484
transform 1 0 21392 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_243
timestamp 1666464484
transform 1 0 28560 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_247
timestamp 1666464484
transform 1 0 29008 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_250
timestamp 1666464484
transform 1 0 29344 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_314
timestamp 1666464484
transform 1 0 36512 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_318
timestamp 1666464484
transform 1 0 36960 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_321
timestamp 1666464484
transform 1 0 37296 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_385
timestamp 1666464484
transform 1 0 44464 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_389
timestamp 1666464484
transform 1 0 44912 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_392
timestamp 1666464484
transform 1 0 45248 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_456
timestamp 1666464484
transform 1 0 52416 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_460
timestamp 1666464484
transform 1 0 52864 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_463
timestamp 1666464484
transform 1 0 53200 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_527
timestamp 1666464484
transform 1 0 60368 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_531
timestamp 1666464484
transform 1 0 60816 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_534
timestamp 1666464484
transform 1 0 61152 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_598
timestamp 1666464484
transform 1 0 68320 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_602
timestamp 1666464484
transform 1 0 68768 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_605
timestamp 1666464484
transform 1 0 69104 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_669
timestamp 1666464484
transform 1 0 76272 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_673
timestamp 1666464484
transform 1 0 76720 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_676
timestamp 1666464484
transform 1 0 77056 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_740
timestamp 1666464484
transform 1 0 84224 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_744
timestamp 1666464484
transform 1 0 84672 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_747
timestamp 1666464484
transform 1 0 85008 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_811
timestamp 1666464484
transform 1 0 92176 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_815
timestamp 1666464484
transform 1 0 92624 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_818
timestamp 1666464484
transform 1 0 92960 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_882
timestamp 1666464484
transform 1 0 100128 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_886
timestamp 1666464484
transform 1 0 100576 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_889
timestamp 1666464484
transform 1 0 100912 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_953
timestamp 1666464484
transform 1 0 108080 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_957
timestamp 1666464484
transform 1 0 108528 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_960
timestamp 1666464484
transform 1 0 108864 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1024
timestamp 1666464484
transform 1 0 116032 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1028
timestamp 1666464484
transform 1 0 116480 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_1031
timestamp 1666464484
transform 1 0 116816 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1095
timestamp 1666464484
transform 1 0 123984 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1099
timestamp 1666464484
transform 1 0 124432 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_1102
timestamp 1666464484
transform 1 0 124768 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1166
timestamp 1666464484
transform 1 0 131936 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1170
timestamp 1666464484
transform 1 0 132384 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_1173
timestamp 1666464484
transform 1 0 132720 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1237
timestamp 1666464484
transform 1 0 139888 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1241
timestamp 1666464484
transform 1 0 140336 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_1244
timestamp 1666464484
transform 1 0 140672 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1308
timestamp 1666464484
transform 1 0 147840 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1312
timestamp 1666464484
transform 1 0 148288 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_1315
timestamp 1666464484
transform 1 0 148624 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1379
timestamp 1666464484
transform 1 0 155792 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1383
timestamp 1666464484
transform 1 0 156240 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_1386
timestamp 1666464484
transform 1 0 156576 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1450
timestamp 1666464484
transform 1 0 163744 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1454
timestamp 1666464484
transform 1 0 164192 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_1457
timestamp 1666464484
transform 1 0 164528 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1521
timestamp 1666464484
transform 1 0 171696 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1525
timestamp 1666464484
transform 1 0 172144 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_102_1528
timestamp 1666464484
transform 1 0 172480 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_1560
timestamp 1666464484
transform 1 0 176064 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1576
timestamp 1666464484
transform 1 0 177856 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1580
timestamp 1666464484
transform 1 0 178304 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_2
timestamp 1666464484
transform 1 0 1568 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_66
timestamp 1666464484
transform 1 0 8736 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_70
timestamp 1666464484
transform 1 0 9184 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_73
timestamp 1666464484
transform 1 0 9520 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_137
timestamp 1666464484
transform 1 0 16688 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_141
timestamp 1666464484
transform 1 0 17136 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_144
timestamp 1666464484
transform 1 0 17472 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_208
timestamp 1666464484
transform 1 0 24640 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_212
timestamp 1666464484
transform 1 0 25088 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_215
timestamp 1666464484
transform 1 0 25424 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_279
timestamp 1666464484
transform 1 0 32592 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_283
timestamp 1666464484
transform 1 0 33040 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_286
timestamp 1666464484
transform 1 0 33376 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_350
timestamp 1666464484
transform 1 0 40544 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_354
timestamp 1666464484
transform 1 0 40992 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_357
timestamp 1666464484
transform 1 0 41328 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_421
timestamp 1666464484
transform 1 0 48496 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_425
timestamp 1666464484
transform 1 0 48944 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_428
timestamp 1666464484
transform 1 0 49280 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_492
timestamp 1666464484
transform 1 0 56448 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_496
timestamp 1666464484
transform 1 0 56896 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_499
timestamp 1666464484
transform 1 0 57232 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_563
timestamp 1666464484
transform 1 0 64400 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_567
timestamp 1666464484
transform 1 0 64848 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_570
timestamp 1666464484
transform 1 0 65184 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_634
timestamp 1666464484
transform 1 0 72352 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_638
timestamp 1666464484
transform 1 0 72800 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_641
timestamp 1666464484
transform 1 0 73136 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_705
timestamp 1666464484
transform 1 0 80304 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_709
timestamp 1666464484
transform 1 0 80752 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_712
timestamp 1666464484
transform 1 0 81088 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_776
timestamp 1666464484
transform 1 0 88256 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_780
timestamp 1666464484
transform 1 0 88704 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_783
timestamp 1666464484
transform 1 0 89040 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_847
timestamp 1666464484
transform 1 0 96208 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_851
timestamp 1666464484
transform 1 0 96656 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_854
timestamp 1666464484
transform 1 0 96992 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_918
timestamp 1666464484
transform 1 0 104160 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_922
timestamp 1666464484
transform 1 0 104608 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_925
timestamp 1666464484
transform 1 0 104944 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_989
timestamp 1666464484
transform 1 0 112112 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_993
timestamp 1666464484
transform 1 0 112560 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_996
timestamp 1666464484
transform 1 0 112896 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1060
timestamp 1666464484
transform 1 0 120064 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1064
timestamp 1666464484
transform 1 0 120512 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_1067
timestamp 1666464484
transform 1 0 120848 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1131
timestamp 1666464484
transform 1 0 128016 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1135
timestamp 1666464484
transform 1 0 128464 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_1138
timestamp 1666464484
transform 1 0 128800 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1202
timestamp 1666464484
transform 1 0 135968 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1206
timestamp 1666464484
transform 1 0 136416 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_1209
timestamp 1666464484
transform 1 0 136752 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1273
timestamp 1666464484
transform 1 0 143920 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1277
timestamp 1666464484
transform 1 0 144368 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_1280
timestamp 1666464484
transform 1 0 144704 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1344
timestamp 1666464484
transform 1 0 151872 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1348
timestamp 1666464484
transform 1 0 152320 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_1351
timestamp 1666464484
transform 1 0 152656 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1415
timestamp 1666464484
transform 1 0 159824 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1419
timestamp 1666464484
transform 1 0 160272 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_1422
timestamp 1666464484
transform 1 0 160608 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1486
timestamp 1666464484
transform 1 0 167776 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1490
timestamp 1666464484
transform 1 0 168224 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_1493
timestamp 1666464484
transform 1 0 168560 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1557
timestamp 1666464484
transform 1 0 175728 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1561
timestamp 1666464484
transform 1 0 176176 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_103_1564
timestamp 1666464484
transform 1 0 176512 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1580
timestamp 1666464484
transform 1 0 178304 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_104_2
timestamp 1666464484
transform 1 0 1568 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_34
timestamp 1666464484
transform 1 0 5152 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_37
timestamp 1666464484
transform 1 0 5488 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_101
timestamp 1666464484
transform 1 0 12656 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_105
timestamp 1666464484
transform 1 0 13104 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_108
timestamp 1666464484
transform 1 0 13440 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_172
timestamp 1666464484
transform 1 0 20608 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_176
timestamp 1666464484
transform 1 0 21056 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_179
timestamp 1666464484
transform 1 0 21392 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_243
timestamp 1666464484
transform 1 0 28560 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_247
timestamp 1666464484
transform 1 0 29008 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_250
timestamp 1666464484
transform 1 0 29344 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_314
timestamp 1666464484
transform 1 0 36512 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_318
timestamp 1666464484
transform 1 0 36960 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_321
timestamp 1666464484
transform 1 0 37296 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_385
timestamp 1666464484
transform 1 0 44464 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_389
timestamp 1666464484
transform 1 0 44912 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_392
timestamp 1666464484
transform 1 0 45248 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_456
timestamp 1666464484
transform 1 0 52416 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_460
timestamp 1666464484
transform 1 0 52864 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_463
timestamp 1666464484
transform 1 0 53200 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_527
timestamp 1666464484
transform 1 0 60368 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_531
timestamp 1666464484
transform 1 0 60816 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_534
timestamp 1666464484
transform 1 0 61152 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_598
timestamp 1666464484
transform 1 0 68320 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_602
timestamp 1666464484
transform 1 0 68768 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_605
timestamp 1666464484
transform 1 0 69104 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_669
timestamp 1666464484
transform 1 0 76272 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_673
timestamp 1666464484
transform 1 0 76720 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_676
timestamp 1666464484
transform 1 0 77056 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_740
timestamp 1666464484
transform 1 0 84224 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_744
timestamp 1666464484
transform 1 0 84672 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_747
timestamp 1666464484
transform 1 0 85008 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_811
timestamp 1666464484
transform 1 0 92176 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_815
timestamp 1666464484
transform 1 0 92624 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_818
timestamp 1666464484
transform 1 0 92960 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_882
timestamp 1666464484
transform 1 0 100128 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_886
timestamp 1666464484
transform 1 0 100576 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_889
timestamp 1666464484
transform 1 0 100912 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_953
timestamp 1666464484
transform 1 0 108080 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_957
timestamp 1666464484
transform 1 0 108528 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_960
timestamp 1666464484
transform 1 0 108864 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1024
timestamp 1666464484
transform 1 0 116032 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1028
timestamp 1666464484
transform 1 0 116480 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_1031
timestamp 1666464484
transform 1 0 116816 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1095
timestamp 1666464484
transform 1 0 123984 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1099
timestamp 1666464484
transform 1 0 124432 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_1102
timestamp 1666464484
transform 1 0 124768 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1166
timestamp 1666464484
transform 1 0 131936 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1170
timestamp 1666464484
transform 1 0 132384 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_1173
timestamp 1666464484
transform 1 0 132720 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1237
timestamp 1666464484
transform 1 0 139888 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1241
timestamp 1666464484
transform 1 0 140336 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_1244
timestamp 1666464484
transform 1 0 140672 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1308
timestamp 1666464484
transform 1 0 147840 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1312
timestamp 1666464484
transform 1 0 148288 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_1315
timestamp 1666464484
transform 1 0 148624 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1379
timestamp 1666464484
transform 1 0 155792 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1383
timestamp 1666464484
transform 1 0 156240 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_1386
timestamp 1666464484
transform 1 0 156576 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1450
timestamp 1666464484
transform 1 0 163744 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1454
timestamp 1666464484
transform 1 0 164192 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_1457
timestamp 1666464484
transform 1 0 164528 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1521
timestamp 1666464484
transform 1 0 171696 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1525
timestamp 1666464484
transform 1 0 172144 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_104_1528
timestamp 1666464484
transform 1 0 172480 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_104_1560
timestamp 1666464484
transform 1 0 176064 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1576
timestamp 1666464484
transform 1 0 177856 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1580
timestamp 1666464484
transform 1 0 178304 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_2
timestamp 1666464484
transform 1 0 1568 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_66
timestamp 1666464484
transform 1 0 8736 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_70
timestamp 1666464484
transform 1 0 9184 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_73
timestamp 1666464484
transform 1 0 9520 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_137
timestamp 1666464484
transform 1 0 16688 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_141
timestamp 1666464484
transform 1 0 17136 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_144
timestamp 1666464484
transform 1 0 17472 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_208
timestamp 1666464484
transform 1 0 24640 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_212
timestamp 1666464484
transform 1 0 25088 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_215
timestamp 1666464484
transform 1 0 25424 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_279
timestamp 1666464484
transform 1 0 32592 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_283
timestamp 1666464484
transform 1 0 33040 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_286
timestamp 1666464484
transform 1 0 33376 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_350
timestamp 1666464484
transform 1 0 40544 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_354
timestamp 1666464484
transform 1 0 40992 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_357
timestamp 1666464484
transform 1 0 41328 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_421
timestamp 1666464484
transform 1 0 48496 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_425
timestamp 1666464484
transform 1 0 48944 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_428
timestamp 1666464484
transform 1 0 49280 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_492
timestamp 1666464484
transform 1 0 56448 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_496
timestamp 1666464484
transform 1 0 56896 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_499
timestamp 1666464484
transform 1 0 57232 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_563
timestamp 1666464484
transform 1 0 64400 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_567
timestamp 1666464484
transform 1 0 64848 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_570
timestamp 1666464484
transform 1 0 65184 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_634
timestamp 1666464484
transform 1 0 72352 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_638
timestamp 1666464484
transform 1 0 72800 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_641
timestamp 1666464484
transform 1 0 73136 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_705
timestamp 1666464484
transform 1 0 80304 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_709
timestamp 1666464484
transform 1 0 80752 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_712
timestamp 1666464484
transform 1 0 81088 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_776
timestamp 1666464484
transform 1 0 88256 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_780
timestamp 1666464484
transform 1 0 88704 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_783
timestamp 1666464484
transform 1 0 89040 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_847
timestamp 1666464484
transform 1 0 96208 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_851
timestamp 1666464484
transform 1 0 96656 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_854
timestamp 1666464484
transform 1 0 96992 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_918
timestamp 1666464484
transform 1 0 104160 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_922
timestamp 1666464484
transform 1 0 104608 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_925
timestamp 1666464484
transform 1 0 104944 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_989
timestamp 1666464484
transform 1 0 112112 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_993
timestamp 1666464484
transform 1 0 112560 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_996
timestamp 1666464484
transform 1 0 112896 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_1060
timestamp 1666464484
transform 1 0 120064 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1064
timestamp 1666464484
transform 1 0 120512 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_1067
timestamp 1666464484
transform 1 0 120848 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_1131
timestamp 1666464484
transform 1 0 128016 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1135
timestamp 1666464484
transform 1 0 128464 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_1138
timestamp 1666464484
transform 1 0 128800 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_1202
timestamp 1666464484
transform 1 0 135968 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1206
timestamp 1666464484
transform 1 0 136416 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_1209
timestamp 1666464484
transform 1 0 136752 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_1273
timestamp 1666464484
transform 1 0 143920 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1277
timestamp 1666464484
transform 1 0 144368 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_1280
timestamp 1666464484
transform 1 0 144704 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_1344
timestamp 1666464484
transform 1 0 151872 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1348
timestamp 1666464484
transform 1 0 152320 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_1351
timestamp 1666464484
transform 1 0 152656 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_1415
timestamp 1666464484
transform 1 0 159824 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1419
timestamp 1666464484
transform 1 0 160272 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_1422
timestamp 1666464484
transform 1 0 160608 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_1486
timestamp 1666464484
transform 1 0 167776 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1490
timestamp 1666464484
transform 1 0 168224 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_1493
timestamp 1666464484
transform 1 0 168560 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_1557
timestamp 1666464484
transform 1 0 175728 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1561
timestamp 1666464484
transform 1 0 176176 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_105_1564
timestamp 1666464484
transform 1 0 176512 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1580
timestamp 1666464484
transform 1 0 178304 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_106_2
timestamp 1666464484
transform 1 0 1568 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_34
timestamp 1666464484
transform 1 0 5152 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_37
timestamp 1666464484
transform 1 0 5488 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_101
timestamp 1666464484
transform 1 0 12656 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_105
timestamp 1666464484
transform 1 0 13104 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_108
timestamp 1666464484
transform 1 0 13440 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_172
timestamp 1666464484
transform 1 0 20608 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_176
timestamp 1666464484
transform 1 0 21056 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_179
timestamp 1666464484
transform 1 0 21392 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_243
timestamp 1666464484
transform 1 0 28560 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_247
timestamp 1666464484
transform 1 0 29008 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_250
timestamp 1666464484
transform 1 0 29344 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_314
timestamp 1666464484
transform 1 0 36512 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_318
timestamp 1666464484
transform 1 0 36960 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_321
timestamp 1666464484
transform 1 0 37296 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_385
timestamp 1666464484
transform 1 0 44464 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_389
timestamp 1666464484
transform 1 0 44912 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_392
timestamp 1666464484
transform 1 0 45248 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_456
timestamp 1666464484
transform 1 0 52416 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_460
timestamp 1666464484
transform 1 0 52864 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_463
timestamp 1666464484
transform 1 0 53200 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_527
timestamp 1666464484
transform 1 0 60368 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_531
timestamp 1666464484
transform 1 0 60816 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_534
timestamp 1666464484
transform 1 0 61152 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_598
timestamp 1666464484
transform 1 0 68320 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_602
timestamp 1666464484
transform 1 0 68768 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_605
timestamp 1666464484
transform 1 0 69104 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_669
timestamp 1666464484
transform 1 0 76272 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_673
timestamp 1666464484
transform 1 0 76720 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_676
timestamp 1666464484
transform 1 0 77056 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_740
timestamp 1666464484
transform 1 0 84224 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_744
timestamp 1666464484
transform 1 0 84672 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_747
timestamp 1666464484
transform 1 0 85008 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_811
timestamp 1666464484
transform 1 0 92176 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_815
timestamp 1666464484
transform 1 0 92624 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_818
timestamp 1666464484
transform 1 0 92960 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_882
timestamp 1666464484
transform 1 0 100128 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_886
timestamp 1666464484
transform 1 0 100576 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_889
timestamp 1666464484
transform 1 0 100912 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_953
timestamp 1666464484
transform 1 0 108080 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_957
timestamp 1666464484
transform 1 0 108528 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_960
timestamp 1666464484
transform 1 0 108864 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1024
timestamp 1666464484
transform 1 0 116032 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1028
timestamp 1666464484
transform 1 0 116480 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_1031
timestamp 1666464484
transform 1 0 116816 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1095
timestamp 1666464484
transform 1 0 123984 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1099
timestamp 1666464484
transform 1 0 124432 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_1102
timestamp 1666464484
transform 1 0 124768 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1166
timestamp 1666464484
transform 1 0 131936 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1170
timestamp 1666464484
transform 1 0 132384 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_1173
timestamp 1666464484
transform 1 0 132720 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1237
timestamp 1666464484
transform 1 0 139888 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1241
timestamp 1666464484
transform 1 0 140336 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_1244
timestamp 1666464484
transform 1 0 140672 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1308
timestamp 1666464484
transform 1 0 147840 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1312
timestamp 1666464484
transform 1 0 148288 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_1315
timestamp 1666464484
transform 1 0 148624 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1379
timestamp 1666464484
transform 1 0 155792 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1383
timestamp 1666464484
transform 1 0 156240 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_1386
timestamp 1666464484
transform 1 0 156576 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1450
timestamp 1666464484
transform 1 0 163744 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1454
timestamp 1666464484
transform 1 0 164192 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_1457
timestamp 1666464484
transform 1 0 164528 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1521
timestamp 1666464484
transform 1 0 171696 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1525
timestamp 1666464484
transform 1 0 172144 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_106_1528
timestamp 1666464484
transform 1 0 172480 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_106_1560
timestamp 1666464484
transform 1 0 176064 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1576
timestamp 1666464484
transform 1 0 177856 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1580
timestamp 1666464484
transform 1 0 178304 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_2
timestamp 1666464484
transform 1 0 1568 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_66
timestamp 1666464484
transform 1 0 8736 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_70
timestamp 1666464484
transform 1 0 9184 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_73
timestamp 1666464484
transform 1 0 9520 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_137
timestamp 1666464484
transform 1 0 16688 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_141
timestamp 1666464484
transform 1 0 17136 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_144
timestamp 1666464484
transform 1 0 17472 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_208
timestamp 1666464484
transform 1 0 24640 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_212
timestamp 1666464484
transform 1 0 25088 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_215
timestamp 1666464484
transform 1 0 25424 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_279
timestamp 1666464484
transform 1 0 32592 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_283
timestamp 1666464484
transform 1 0 33040 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_286
timestamp 1666464484
transform 1 0 33376 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_350
timestamp 1666464484
transform 1 0 40544 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_354
timestamp 1666464484
transform 1 0 40992 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_357
timestamp 1666464484
transform 1 0 41328 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_421
timestamp 1666464484
transform 1 0 48496 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_425
timestamp 1666464484
transform 1 0 48944 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_428
timestamp 1666464484
transform 1 0 49280 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_492
timestamp 1666464484
transform 1 0 56448 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_496
timestamp 1666464484
transform 1 0 56896 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_499
timestamp 1666464484
transform 1 0 57232 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_563
timestamp 1666464484
transform 1 0 64400 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_567
timestamp 1666464484
transform 1 0 64848 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_570
timestamp 1666464484
transform 1 0 65184 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_634
timestamp 1666464484
transform 1 0 72352 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_638
timestamp 1666464484
transform 1 0 72800 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_641
timestamp 1666464484
transform 1 0 73136 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_705
timestamp 1666464484
transform 1 0 80304 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_709
timestamp 1666464484
transform 1 0 80752 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_712
timestamp 1666464484
transform 1 0 81088 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_776
timestamp 1666464484
transform 1 0 88256 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_780
timestamp 1666464484
transform 1 0 88704 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_783
timestamp 1666464484
transform 1 0 89040 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_847
timestamp 1666464484
transform 1 0 96208 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_851
timestamp 1666464484
transform 1 0 96656 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_854
timestamp 1666464484
transform 1 0 96992 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_918
timestamp 1666464484
transform 1 0 104160 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_922
timestamp 1666464484
transform 1 0 104608 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_925
timestamp 1666464484
transform 1 0 104944 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_989
timestamp 1666464484
transform 1 0 112112 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_993
timestamp 1666464484
transform 1 0 112560 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_996
timestamp 1666464484
transform 1 0 112896 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1060
timestamp 1666464484
transform 1 0 120064 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1064
timestamp 1666464484
transform 1 0 120512 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_1067
timestamp 1666464484
transform 1 0 120848 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1131
timestamp 1666464484
transform 1 0 128016 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1135
timestamp 1666464484
transform 1 0 128464 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_1138
timestamp 1666464484
transform 1 0 128800 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1202
timestamp 1666464484
transform 1 0 135968 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1206
timestamp 1666464484
transform 1 0 136416 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_1209
timestamp 1666464484
transform 1 0 136752 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1273
timestamp 1666464484
transform 1 0 143920 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1277
timestamp 1666464484
transform 1 0 144368 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_1280
timestamp 1666464484
transform 1 0 144704 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1344
timestamp 1666464484
transform 1 0 151872 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1348
timestamp 1666464484
transform 1 0 152320 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_1351
timestamp 1666464484
transform 1 0 152656 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1415
timestamp 1666464484
transform 1 0 159824 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1419
timestamp 1666464484
transform 1 0 160272 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_1422
timestamp 1666464484
transform 1 0 160608 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1486
timestamp 1666464484
transform 1 0 167776 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1490
timestamp 1666464484
transform 1 0 168224 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_1493
timestamp 1666464484
transform 1 0 168560 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_1557
timestamp 1666464484
transform 1 0 175728 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1561
timestamp 1666464484
transform 1 0 176176 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_107_1564
timestamp 1666464484
transform 1 0 176512 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1580
timestamp 1666464484
transform 1 0 178304 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_108_2
timestamp 1666464484
transform 1 0 1568 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_34
timestamp 1666464484
transform 1 0 5152 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_37
timestamp 1666464484
transform 1 0 5488 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_101
timestamp 1666464484
transform 1 0 12656 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_105
timestamp 1666464484
transform 1 0 13104 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_108
timestamp 1666464484
transform 1 0 13440 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_172
timestamp 1666464484
transform 1 0 20608 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_176
timestamp 1666464484
transform 1 0 21056 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_179
timestamp 1666464484
transform 1 0 21392 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_243
timestamp 1666464484
transform 1 0 28560 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_247
timestamp 1666464484
transform 1 0 29008 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_250
timestamp 1666464484
transform 1 0 29344 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_314
timestamp 1666464484
transform 1 0 36512 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_318
timestamp 1666464484
transform 1 0 36960 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_321
timestamp 1666464484
transform 1 0 37296 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_385
timestamp 1666464484
transform 1 0 44464 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_389
timestamp 1666464484
transform 1 0 44912 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_392
timestamp 1666464484
transform 1 0 45248 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_456
timestamp 1666464484
transform 1 0 52416 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_460
timestamp 1666464484
transform 1 0 52864 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_463
timestamp 1666464484
transform 1 0 53200 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_527
timestamp 1666464484
transform 1 0 60368 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_531
timestamp 1666464484
transform 1 0 60816 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_534
timestamp 1666464484
transform 1 0 61152 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_598
timestamp 1666464484
transform 1 0 68320 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_602
timestamp 1666464484
transform 1 0 68768 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_605
timestamp 1666464484
transform 1 0 69104 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_669
timestamp 1666464484
transform 1 0 76272 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_673
timestamp 1666464484
transform 1 0 76720 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_676
timestamp 1666464484
transform 1 0 77056 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_740
timestamp 1666464484
transform 1 0 84224 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_744
timestamp 1666464484
transform 1 0 84672 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_747
timestamp 1666464484
transform 1 0 85008 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_811
timestamp 1666464484
transform 1 0 92176 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_815
timestamp 1666464484
transform 1 0 92624 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_818
timestamp 1666464484
transform 1 0 92960 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_882
timestamp 1666464484
transform 1 0 100128 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_886
timestamp 1666464484
transform 1 0 100576 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_889
timestamp 1666464484
transform 1 0 100912 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_953
timestamp 1666464484
transform 1 0 108080 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_957
timestamp 1666464484
transform 1 0 108528 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_960
timestamp 1666464484
transform 1 0 108864 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1024
timestamp 1666464484
transform 1 0 116032 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1028
timestamp 1666464484
transform 1 0 116480 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_1031
timestamp 1666464484
transform 1 0 116816 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1095
timestamp 1666464484
transform 1 0 123984 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1099
timestamp 1666464484
transform 1 0 124432 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_1102
timestamp 1666464484
transform 1 0 124768 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1166
timestamp 1666464484
transform 1 0 131936 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1170
timestamp 1666464484
transform 1 0 132384 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_1173
timestamp 1666464484
transform 1 0 132720 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1237
timestamp 1666464484
transform 1 0 139888 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1241
timestamp 1666464484
transform 1 0 140336 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_1244
timestamp 1666464484
transform 1 0 140672 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1308
timestamp 1666464484
transform 1 0 147840 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1312
timestamp 1666464484
transform 1 0 148288 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_1315
timestamp 1666464484
transform 1 0 148624 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1379
timestamp 1666464484
transform 1 0 155792 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1383
timestamp 1666464484
transform 1 0 156240 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_1386
timestamp 1666464484
transform 1 0 156576 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1450
timestamp 1666464484
transform 1 0 163744 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1454
timestamp 1666464484
transform 1 0 164192 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_1457
timestamp 1666464484
transform 1 0 164528 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1521
timestamp 1666464484
transform 1 0 171696 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1525
timestamp 1666464484
transform 1 0 172144 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_108_1528
timestamp 1666464484
transform 1 0 172480 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_108_1560
timestamp 1666464484
transform 1 0 176064 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1576
timestamp 1666464484
transform 1 0 177856 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1580
timestamp 1666464484
transform 1 0 178304 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_2
timestamp 1666464484
transform 1 0 1568 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_66
timestamp 1666464484
transform 1 0 8736 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_70
timestamp 1666464484
transform 1 0 9184 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_73
timestamp 1666464484
transform 1 0 9520 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_137
timestamp 1666464484
transform 1 0 16688 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_141
timestamp 1666464484
transform 1 0 17136 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_144
timestamp 1666464484
transform 1 0 17472 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_208
timestamp 1666464484
transform 1 0 24640 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_212
timestamp 1666464484
transform 1 0 25088 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_215
timestamp 1666464484
transform 1 0 25424 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_279
timestamp 1666464484
transform 1 0 32592 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_283
timestamp 1666464484
transform 1 0 33040 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_286
timestamp 1666464484
transform 1 0 33376 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_350
timestamp 1666464484
transform 1 0 40544 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_354
timestamp 1666464484
transform 1 0 40992 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_357
timestamp 1666464484
transform 1 0 41328 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_421
timestamp 1666464484
transform 1 0 48496 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_425
timestamp 1666464484
transform 1 0 48944 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_428
timestamp 1666464484
transform 1 0 49280 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_492
timestamp 1666464484
transform 1 0 56448 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_496
timestamp 1666464484
transform 1 0 56896 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_499
timestamp 1666464484
transform 1 0 57232 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_563
timestamp 1666464484
transform 1 0 64400 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_567
timestamp 1666464484
transform 1 0 64848 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_570
timestamp 1666464484
transform 1 0 65184 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_634
timestamp 1666464484
transform 1 0 72352 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_638
timestamp 1666464484
transform 1 0 72800 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_641
timestamp 1666464484
transform 1 0 73136 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_705
timestamp 1666464484
transform 1 0 80304 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_709
timestamp 1666464484
transform 1 0 80752 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_712
timestamp 1666464484
transform 1 0 81088 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_776
timestamp 1666464484
transform 1 0 88256 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_780
timestamp 1666464484
transform 1 0 88704 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_783
timestamp 1666464484
transform 1 0 89040 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_847
timestamp 1666464484
transform 1 0 96208 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_851
timestamp 1666464484
transform 1 0 96656 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_854
timestamp 1666464484
transform 1 0 96992 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_918
timestamp 1666464484
transform 1 0 104160 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_922
timestamp 1666464484
transform 1 0 104608 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_925
timestamp 1666464484
transform 1 0 104944 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_989
timestamp 1666464484
transform 1 0 112112 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_993
timestamp 1666464484
transform 1 0 112560 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_996
timestamp 1666464484
transform 1 0 112896 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_1060
timestamp 1666464484
transform 1 0 120064 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1064
timestamp 1666464484
transform 1 0 120512 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_1067
timestamp 1666464484
transform 1 0 120848 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_1131
timestamp 1666464484
transform 1 0 128016 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1135
timestamp 1666464484
transform 1 0 128464 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_1138
timestamp 1666464484
transform 1 0 128800 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_1202
timestamp 1666464484
transform 1 0 135968 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1206
timestamp 1666464484
transform 1 0 136416 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_1209
timestamp 1666464484
transform 1 0 136752 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_1273
timestamp 1666464484
transform 1 0 143920 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1277
timestamp 1666464484
transform 1 0 144368 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_1280
timestamp 1666464484
transform 1 0 144704 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_1344
timestamp 1666464484
transform 1 0 151872 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1348
timestamp 1666464484
transform 1 0 152320 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_1351
timestamp 1666464484
transform 1 0 152656 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_1415
timestamp 1666464484
transform 1 0 159824 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1419
timestamp 1666464484
transform 1 0 160272 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_1422
timestamp 1666464484
transform 1 0 160608 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_1486
timestamp 1666464484
transform 1 0 167776 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1490
timestamp 1666464484
transform 1 0 168224 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_1493
timestamp 1666464484
transform 1 0 168560 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_1557
timestamp 1666464484
transform 1 0 175728 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1561
timestamp 1666464484
transform 1 0 176176 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_1564
timestamp 1666464484
transform 1 0 176512 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1580
timestamp 1666464484
transform 1 0 178304 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_110_2
timestamp 1666464484
transform 1 0 1568 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_34
timestamp 1666464484
transform 1 0 5152 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_37
timestamp 1666464484
transform 1 0 5488 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_101
timestamp 1666464484
transform 1 0 12656 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_105
timestamp 1666464484
transform 1 0 13104 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_108
timestamp 1666464484
transform 1 0 13440 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_172
timestamp 1666464484
transform 1 0 20608 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_176
timestamp 1666464484
transform 1 0 21056 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_179
timestamp 1666464484
transform 1 0 21392 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_243
timestamp 1666464484
transform 1 0 28560 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_247
timestamp 1666464484
transform 1 0 29008 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_250
timestamp 1666464484
transform 1 0 29344 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_314
timestamp 1666464484
transform 1 0 36512 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_318
timestamp 1666464484
transform 1 0 36960 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_321
timestamp 1666464484
transform 1 0 37296 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_385
timestamp 1666464484
transform 1 0 44464 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_389
timestamp 1666464484
transform 1 0 44912 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_392
timestamp 1666464484
transform 1 0 45248 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_456
timestamp 1666464484
transform 1 0 52416 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_460
timestamp 1666464484
transform 1 0 52864 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_463
timestamp 1666464484
transform 1 0 53200 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_527
timestamp 1666464484
transform 1 0 60368 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_531
timestamp 1666464484
transform 1 0 60816 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_534
timestamp 1666464484
transform 1 0 61152 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_598
timestamp 1666464484
transform 1 0 68320 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_602
timestamp 1666464484
transform 1 0 68768 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_605
timestamp 1666464484
transform 1 0 69104 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_669
timestamp 1666464484
transform 1 0 76272 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_673
timestamp 1666464484
transform 1 0 76720 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_676
timestamp 1666464484
transform 1 0 77056 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_740
timestamp 1666464484
transform 1 0 84224 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_744
timestamp 1666464484
transform 1 0 84672 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_747
timestamp 1666464484
transform 1 0 85008 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_811
timestamp 1666464484
transform 1 0 92176 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_815
timestamp 1666464484
transform 1 0 92624 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_818
timestamp 1666464484
transform 1 0 92960 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_882
timestamp 1666464484
transform 1 0 100128 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_886
timestamp 1666464484
transform 1 0 100576 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_889
timestamp 1666464484
transform 1 0 100912 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_953
timestamp 1666464484
transform 1 0 108080 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_957
timestamp 1666464484
transform 1 0 108528 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_960
timestamp 1666464484
transform 1 0 108864 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1024
timestamp 1666464484
transform 1 0 116032 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1028
timestamp 1666464484
transform 1 0 116480 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_1031
timestamp 1666464484
transform 1 0 116816 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1095
timestamp 1666464484
transform 1 0 123984 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1099
timestamp 1666464484
transform 1 0 124432 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_1102
timestamp 1666464484
transform 1 0 124768 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1166
timestamp 1666464484
transform 1 0 131936 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1170
timestamp 1666464484
transform 1 0 132384 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_1173
timestamp 1666464484
transform 1 0 132720 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1237
timestamp 1666464484
transform 1 0 139888 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1241
timestamp 1666464484
transform 1 0 140336 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_1244
timestamp 1666464484
transform 1 0 140672 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1308
timestamp 1666464484
transform 1 0 147840 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1312
timestamp 1666464484
transform 1 0 148288 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_1315
timestamp 1666464484
transform 1 0 148624 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1379
timestamp 1666464484
transform 1 0 155792 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1383
timestamp 1666464484
transform 1 0 156240 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_1386
timestamp 1666464484
transform 1 0 156576 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1450
timestamp 1666464484
transform 1 0 163744 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1454
timestamp 1666464484
transform 1 0 164192 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_1457
timestamp 1666464484
transform 1 0 164528 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1521
timestamp 1666464484
transform 1 0 171696 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1525
timestamp 1666464484
transform 1 0 172144 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_110_1528
timestamp 1666464484
transform 1 0 172480 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_110_1560
timestamp 1666464484
transform 1 0 176064 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1576
timestamp 1666464484
transform 1 0 177856 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1580
timestamp 1666464484
transform 1 0 178304 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_2
timestamp 1666464484
transform 1 0 1568 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_66
timestamp 1666464484
transform 1 0 8736 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_70
timestamp 1666464484
transform 1 0 9184 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_73
timestamp 1666464484
transform 1 0 9520 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_137
timestamp 1666464484
transform 1 0 16688 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_141
timestamp 1666464484
transform 1 0 17136 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_144
timestamp 1666464484
transform 1 0 17472 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_208
timestamp 1666464484
transform 1 0 24640 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_212
timestamp 1666464484
transform 1 0 25088 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_215
timestamp 1666464484
transform 1 0 25424 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_279
timestamp 1666464484
transform 1 0 32592 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_283
timestamp 1666464484
transform 1 0 33040 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_286
timestamp 1666464484
transform 1 0 33376 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_350
timestamp 1666464484
transform 1 0 40544 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_354
timestamp 1666464484
transform 1 0 40992 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_357
timestamp 1666464484
transform 1 0 41328 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_421
timestamp 1666464484
transform 1 0 48496 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_425
timestamp 1666464484
transform 1 0 48944 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_428
timestamp 1666464484
transform 1 0 49280 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_492
timestamp 1666464484
transform 1 0 56448 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_496
timestamp 1666464484
transform 1 0 56896 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_499
timestamp 1666464484
transform 1 0 57232 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_563
timestamp 1666464484
transform 1 0 64400 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_567
timestamp 1666464484
transform 1 0 64848 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_570
timestamp 1666464484
transform 1 0 65184 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_634
timestamp 1666464484
transform 1 0 72352 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_638
timestamp 1666464484
transform 1 0 72800 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_641
timestamp 1666464484
transform 1 0 73136 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_705
timestamp 1666464484
transform 1 0 80304 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_709
timestamp 1666464484
transform 1 0 80752 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_712
timestamp 1666464484
transform 1 0 81088 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_776
timestamp 1666464484
transform 1 0 88256 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_780
timestamp 1666464484
transform 1 0 88704 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_783
timestamp 1666464484
transform 1 0 89040 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_847
timestamp 1666464484
transform 1 0 96208 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_851
timestamp 1666464484
transform 1 0 96656 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_854
timestamp 1666464484
transform 1 0 96992 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_918
timestamp 1666464484
transform 1 0 104160 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_922
timestamp 1666464484
transform 1 0 104608 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_925
timestamp 1666464484
transform 1 0 104944 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_989
timestamp 1666464484
transform 1 0 112112 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_993
timestamp 1666464484
transform 1 0 112560 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_996
timestamp 1666464484
transform 1 0 112896 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_1060
timestamp 1666464484
transform 1 0 120064 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1064
timestamp 1666464484
transform 1 0 120512 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_1067
timestamp 1666464484
transform 1 0 120848 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_1131
timestamp 1666464484
transform 1 0 128016 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1135
timestamp 1666464484
transform 1 0 128464 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_1138
timestamp 1666464484
transform 1 0 128800 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_1202
timestamp 1666464484
transform 1 0 135968 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1206
timestamp 1666464484
transform 1 0 136416 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_1209
timestamp 1666464484
transform 1 0 136752 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_1273
timestamp 1666464484
transform 1 0 143920 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1277
timestamp 1666464484
transform 1 0 144368 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_1280
timestamp 1666464484
transform 1 0 144704 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_1344
timestamp 1666464484
transform 1 0 151872 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1348
timestamp 1666464484
transform 1 0 152320 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_1351
timestamp 1666464484
transform 1 0 152656 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_1415
timestamp 1666464484
transform 1 0 159824 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1419
timestamp 1666464484
transform 1 0 160272 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_1422
timestamp 1666464484
transform 1 0 160608 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_1486
timestamp 1666464484
transform 1 0 167776 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1490
timestamp 1666464484
transform 1 0 168224 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_1493
timestamp 1666464484
transform 1 0 168560 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_1557
timestamp 1666464484
transform 1 0 175728 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1561
timestamp 1666464484
transform 1 0 176176 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_111_1564
timestamp 1666464484
transform 1 0 176512 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1580
timestamp 1666464484
transform 1 0 178304 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_112_2
timestamp 1666464484
transform 1 0 1568 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_34
timestamp 1666464484
transform 1 0 5152 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_37
timestamp 1666464484
transform 1 0 5488 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_101
timestamp 1666464484
transform 1 0 12656 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_105
timestamp 1666464484
transform 1 0 13104 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_108
timestamp 1666464484
transform 1 0 13440 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_172
timestamp 1666464484
transform 1 0 20608 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_176
timestamp 1666464484
transform 1 0 21056 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_179
timestamp 1666464484
transform 1 0 21392 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_243
timestamp 1666464484
transform 1 0 28560 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_247
timestamp 1666464484
transform 1 0 29008 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_250
timestamp 1666464484
transform 1 0 29344 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_314
timestamp 1666464484
transform 1 0 36512 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_318
timestamp 1666464484
transform 1 0 36960 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_321
timestamp 1666464484
transform 1 0 37296 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_385
timestamp 1666464484
transform 1 0 44464 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_389
timestamp 1666464484
transform 1 0 44912 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_392
timestamp 1666464484
transform 1 0 45248 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_456
timestamp 1666464484
transform 1 0 52416 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_460
timestamp 1666464484
transform 1 0 52864 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_463
timestamp 1666464484
transform 1 0 53200 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_527
timestamp 1666464484
transform 1 0 60368 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_531
timestamp 1666464484
transform 1 0 60816 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_534
timestamp 1666464484
transform 1 0 61152 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_598
timestamp 1666464484
transform 1 0 68320 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_602
timestamp 1666464484
transform 1 0 68768 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_605
timestamp 1666464484
transform 1 0 69104 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_669
timestamp 1666464484
transform 1 0 76272 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_673
timestamp 1666464484
transform 1 0 76720 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_676
timestamp 1666464484
transform 1 0 77056 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_740
timestamp 1666464484
transform 1 0 84224 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_744
timestamp 1666464484
transform 1 0 84672 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_747
timestamp 1666464484
transform 1 0 85008 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_811
timestamp 1666464484
transform 1 0 92176 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_815
timestamp 1666464484
transform 1 0 92624 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_818
timestamp 1666464484
transform 1 0 92960 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_882
timestamp 1666464484
transform 1 0 100128 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_886
timestamp 1666464484
transform 1 0 100576 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_889
timestamp 1666464484
transform 1 0 100912 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_953
timestamp 1666464484
transform 1 0 108080 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_957
timestamp 1666464484
transform 1 0 108528 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_960
timestamp 1666464484
transform 1 0 108864 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1024
timestamp 1666464484
transform 1 0 116032 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1028
timestamp 1666464484
transform 1 0 116480 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_1031
timestamp 1666464484
transform 1 0 116816 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1095
timestamp 1666464484
transform 1 0 123984 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1099
timestamp 1666464484
transform 1 0 124432 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_1102
timestamp 1666464484
transform 1 0 124768 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1166
timestamp 1666464484
transform 1 0 131936 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1170
timestamp 1666464484
transform 1 0 132384 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_1173
timestamp 1666464484
transform 1 0 132720 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1237
timestamp 1666464484
transform 1 0 139888 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1241
timestamp 1666464484
transform 1 0 140336 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_1244
timestamp 1666464484
transform 1 0 140672 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1308
timestamp 1666464484
transform 1 0 147840 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1312
timestamp 1666464484
transform 1 0 148288 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_1315
timestamp 1666464484
transform 1 0 148624 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1379
timestamp 1666464484
transform 1 0 155792 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1383
timestamp 1666464484
transform 1 0 156240 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_1386
timestamp 1666464484
transform 1 0 156576 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1450
timestamp 1666464484
transform 1 0 163744 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1454
timestamp 1666464484
transform 1 0 164192 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_1457
timestamp 1666464484
transform 1 0 164528 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1521
timestamp 1666464484
transform 1 0 171696 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1525
timestamp 1666464484
transform 1 0 172144 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_112_1528
timestamp 1666464484
transform 1 0 172480 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_112_1560
timestamp 1666464484
transform 1 0 176064 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1576
timestamp 1666464484
transform 1 0 177856 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1580
timestamp 1666464484
transform 1 0 178304 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_2
timestamp 1666464484
transform 1 0 1568 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_66
timestamp 1666464484
transform 1 0 8736 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_70
timestamp 1666464484
transform 1 0 9184 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_73
timestamp 1666464484
transform 1 0 9520 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_137
timestamp 1666464484
transform 1 0 16688 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_141
timestamp 1666464484
transform 1 0 17136 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_144
timestamp 1666464484
transform 1 0 17472 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_208
timestamp 1666464484
transform 1 0 24640 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_212
timestamp 1666464484
transform 1 0 25088 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_215
timestamp 1666464484
transform 1 0 25424 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_279
timestamp 1666464484
transform 1 0 32592 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_283
timestamp 1666464484
transform 1 0 33040 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_286
timestamp 1666464484
transform 1 0 33376 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_350
timestamp 1666464484
transform 1 0 40544 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_354
timestamp 1666464484
transform 1 0 40992 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_357
timestamp 1666464484
transform 1 0 41328 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_421
timestamp 1666464484
transform 1 0 48496 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_425
timestamp 1666464484
transform 1 0 48944 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_428
timestamp 1666464484
transform 1 0 49280 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_492
timestamp 1666464484
transform 1 0 56448 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_496
timestamp 1666464484
transform 1 0 56896 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_499
timestamp 1666464484
transform 1 0 57232 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_563
timestamp 1666464484
transform 1 0 64400 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_567
timestamp 1666464484
transform 1 0 64848 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_570
timestamp 1666464484
transform 1 0 65184 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_634
timestamp 1666464484
transform 1 0 72352 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_638
timestamp 1666464484
transform 1 0 72800 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_641
timestamp 1666464484
transform 1 0 73136 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_705
timestamp 1666464484
transform 1 0 80304 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_709
timestamp 1666464484
transform 1 0 80752 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_712
timestamp 1666464484
transform 1 0 81088 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_776
timestamp 1666464484
transform 1 0 88256 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_780
timestamp 1666464484
transform 1 0 88704 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_783
timestamp 1666464484
transform 1 0 89040 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_847
timestamp 1666464484
transform 1 0 96208 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_851
timestamp 1666464484
transform 1 0 96656 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_854
timestamp 1666464484
transform 1 0 96992 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_918
timestamp 1666464484
transform 1 0 104160 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_922
timestamp 1666464484
transform 1 0 104608 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_925
timestamp 1666464484
transform 1 0 104944 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_989
timestamp 1666464484
transform 1 0 112112 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_993
timestamp 1666464484
transform 1 0 112560 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_996
timestamp 1666464484
transform 1 0 112896 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_1060
timestamp 1666464484
transform 1 0 120064 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1064
timestamp 1666464484
transform 1 0 120512 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_1067
timestamp 1666464484
transform 1 0 120848 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_1131
timestamp 1666464484
transform 1 0 128016 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1135
timestamp 1666464484
transform 1 0 128464 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_1138
timestamp 1666464484
transform 1 0 128800 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_1202
timestamp 1666464484
transform 1 0 135968 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1206
timestamp 1666464484
transform 1 0 136416 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_1209
timestamp 1666464484
transform 1 0 136752 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_1273
timestamp 1666464484
transform 1 0 143920 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1277
timestamp 1666464484
transform 1 0 144368 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_1280
timestamp 1666464484
transform 1 0 144704 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_1344
timestamp 1666464484
transform 1 0 151872 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1348
timestamp 1666464484
transform 1 0 152320 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_1351
timestamp 1666464484
transform 1 0 152656 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_1415
timestamp 1666464484
transform 1 0 159824 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1419
timestamp 1666464484
transform 1 0 160272 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_1422
timestamp 1666464484
transform 1 0 160608 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_1486
timestamp 1666464484
transform 1 0 167776 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1490
timestamp 1666464484
transform 1 0 168224 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_1493
timestamp 1666464484
transform 1 0 168560 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_1557
timestamp 1666464484
transform 1 0 175728 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1561
timestamp 1666464484
transform 1 0 176176 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_113_1564
timestamp 1666464484
transform 1 0 176512 0 -1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1580
timestamp 1666464484
transform 1 0 178304 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_114_2
timestamp 1666464484
transform 1 0 1568 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_34
timestamp 1666464484
transform 1 0 5152 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_37
timestamp 1666464484
transform 1 0 5488 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_101
timestamp 1666464484
transform 1 0 12656 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_105
timestamp 1666464484
transform 1 0 13104 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_108
timestamp 1666464484
transform 1 0 13440 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_172
timestamp 1666464484
transform 1 0 20608 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_176
timestamp 1666464484
transform 1 0 21056 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_179
timestamp 1666464484
transform 1 0 21392 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_243
timestamp 1666464484
transform 1 0 28560 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_247
timestamp 1666464484
transform 1 0 29008 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_250
timestamp 1666464484
transform 1 0 29344 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_314
timestamp 1666464484
transform 1 0 36512 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_318
timestamp 1666464484
transform 1 0 36960 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_321
timestamp 1666464484
transform 1 0 37296 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_385
timestamp 1666464484
transform 1 0 44464 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_389
timestamp 1666464484
transform 1 0 44912 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_392
timestamp 1666464484
transform 1 0 45248 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_456
timestamp 1666464484
transform 1 0 52416 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_460
timestamp 1666464484
transform 1 0 52864 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_463
timestamp 1666464484
transform 1 0 53200 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_527
timestamp 1666464484
transform 1 0 60368 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_531
timestamp 1666464484
transform 1 0 60816 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_534
timestamp 1666464484
transform 1 0 61152 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_598
timestamp 1666464484
transform 1 0 68320 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_602
timestamp 1666464484
transform 1 0 68768 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_605
timestamp 1666464484
transform 1 0 69104 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_669
timestamp 1666464484
transform 1 0 76272 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_673
timestamp 1666464484
transform 1 0 76720 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_676
timestamp 1666464484
transform 1 0 77056 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_740
timestamp 1666464484
transform 1 0 84224 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_744
timestamp 1666464484
transform 1 0 84672 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_747
timestamp 1666464484
transform 1 0 85008 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_811
timestamp 1666464484
transform 1 0 92176 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_815
timestamp 1666464484
transform 1 0 92624 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_818
timestamp 1666464484
transform 1 0 92960 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_882
timestamp 1666464484
transform 1 0 100128 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_886
timestamp 1666464484
transform 1 0 100576 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_889
timestamp 1666464484
transform 1 0 100912 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_953
timestamp 1666464484
transform 1 0 108080 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_957
timestamp 1666464484
transform 1 0 108528 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_960
timestamp 1666464484
transform 1 0 108864 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1024
timestamp 1666464484
transform 1 0 116032 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1028
timestamp 1666464484
transform 1 0 116480 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_1031
timestamp 1666464484
transform 1 0 116816 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1095
timestamp 1666464484
transform 1 0 123984 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1099
timestamp 1666464484
transform 1 0 124432 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_1102
timestamp 1666464484
transform 1 0 124768 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1166
timestamp 1666464484
transform 1 0 131936 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1170
timestamp 1666464484
transform 1 0 132384 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_1173
timestamp 1666464484
transform 1 0 132720 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1237
timestamp 1666464484
transform 1 0 139888 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1241
timestamp 1666464484
transform 1 0 140336 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_1244
timestamp 1666464484
transform 1 0 140672 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1308
timestamp 1666464484
transform 1 0 147840 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1312
timestamp 1666464484
transform 1 0 148288 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_1315
timestamp 1666464484
transform 1 0 148624 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1379
timestamp 1666464484
transform 1 0 155792 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1383
timestamp 1666464484
transform 1 0 156240 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_1386
timestamp 1666464484
transform 1 0 156576 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1450
timestamp 1666464484
transform 1 0 163744 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1454
timestamp 1666464484
transform 1 0 164192 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_1457
timestamp 1666464484
transform 1 0 164528 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1521
timestamp 1666464484
transform 1 0 171696 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1525
timestamp 1666464484
transform 1 0 172144 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_114_1528
timestamp 1666464484
transform 1 0 172480 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_114_1560
timestamp 1666464484
transform 1 0 176064 0 1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1576
timestamp 1666464484
transform 1 0 177856 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1580
timestamp 1666464484
transform 1 0 178304 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_2
timestamp 1666464484
transform 1 0 1568 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_66
timestamp 1666464484
transform 1 0 8736 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_70
timestamp 1666464484
transform 1 0 9184 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_73
timestamp 1666464484
transform 1 0 9520 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_137
timestamp 1666464484
transform 1 0 16688 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_141
timestamp 1666464484
transform 1 0 17136 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_144
timestamp 1666464484
transform 1 0 17472 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_208
timestamp 1666464484
transform 1 0 24640 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_212
timestamp 1666464484
transform 1 0 25088 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_215
timestamp 1666464484
transform 1 0 25424 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_279
timestamp 1666464484
transform 1 0 32592 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_283
timestamp 1666464484
transform 1 0 33040 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_286
timestamp 1666464484
transform 1 0 33376 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_350
timestamp 1666464484
transform 1 0 40544 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_354
timestamp 1666464484
transform 1 0 40992 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_357
timestamp 1666464484
transform 1 0 41328 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_421
timestamp 1666464484
transform 1 0 48496 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_425
timestamp 1666464484
transform 1 0 48944 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_428
timestamp 1666464484
transform 1 0 49280 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_492
timestamp 1666464484
transform 1 0 56448 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_496
timestamp 1666464484
transform 1 0 56896 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_499
timestamp 1666464484
transform 1 0 57232 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_563
timestamp 1666464484
transform 1 0 64400 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_567
timestamp 1666464484
transform 1 0 64848 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_570
timestamp 1666464484
transform 1 0 65184 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_634
timestamp 1666464484
transform 1 0 72352 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_638
timestamp 1666464484
transform 1 0 72800 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_641
timestamp 1666464484
transform 1 0 73136 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_705
timestamp 1666464484
transform 1 0 80304 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_709
timestamp 1666464484
transform 1 0 80752 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_712
timestamp 1666464484
transform 1 0 81088 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_776
timestamp 1666464484
transform 1 0 88256 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_780
timestamp 1666464484
transform 1 0 88704 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_783
timestamp 1666464484
transform 1 0 89040 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_847
timestamp 1666464484
transform 1 0 96208 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_851
timestamp 1666464484
transform 1 0 96656 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_854
timestamp 1666464484
transform 1 0 96992 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_918
timestamp 1666464484
transform 1 0 104160 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_922
timestamp 1666464484
transform 1 0 104608 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_925
timestamp 1666464484
transform 1 0 104944 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_989
timestamp 1666464484
transform 1 0 112112 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_993
timestamp 1666464484
transform 1 0 112560 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_996
timestamp 1666464484
transform 1 0 112896 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_1060
timestamp 1666464484
transform 1 0 120064 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1064
timestamp 1666464484
transform 1 0 120512 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_1067
timestamp 1666464484
transform 1 0 120848 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_1131
timestamp 1666464484
transform 1 0 128016 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1135
timestamp 1666464484
transform 1 0 128464 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_1138
timestamp 1666464484
transform 1 0 128800 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_1202
timestamp 1666464484
transform 1 0 135968 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1206
timestamp 1666464484
transform 1 0 136416 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_1209
timestamp 1666464484
transform 1 0 136752 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_1273
timestamp 1666464484
transform 1 0 143920 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1277
timestamp 1666464484
transform 1 0 144368 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_1280
timestamp 1666464484
transform 1 0 144704 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_1344
timestamp 1666464484
transform 1 0 151872 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1348
timestamp 1666464484
transform 1 0 152320 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_1351
timestamp 1666464484
transform 1 0 152656 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_1415
timestamp 1666464484
transform 1 0 159824 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1419
timestamp 1666464484
transform 1 0 160272 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_1422
timestamp 1666464484
transform 1 0 160608 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_1486
timestamp 1666464484
transform 1 0 167776 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1490
timestamp 1666464484
transform 1 0 168224 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_1493
timestamp 1666464484
transform 1 0 168560 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_1557
timestamp 1666464484
transform 1 0 175728 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1561
timestamp 1666464484
transform 1 0 176176 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_115_1564
timestamp 1666464484
transform 1 0 176512 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1580
timestamp 1666464484
transform 1 0 178304 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_116_2
timestamp 1666464484
transform 1 0 1568 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_34
timestamp 1666464484
transform 1 0 5152 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_37
timestamp 1666464484
transform 1 0 5488 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_101
timestamp 1666464484
transform 1 0 12656 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_105
timestamp 1666464484
transform 1 0 13104 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_108
timestamp 1666464484
transform 1 0 13440 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_172
timestamp 1666464484
transform 1 0 20608 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_176
timestamp 1666464484
transform 1 0 21056 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_179
timestamp 1666464484
transform 1 0 21392 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_243
timestamp 1666464484
transform 1 0 28560 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_247
timestamp 1666464484
transform 1 0 29008 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_250
timestamp 1666464484
transform 1 0 29344 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_314
timestamp 1666464484
transform 1 0 36512 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_318
timestamp 1666464484
transform 1 0 36960 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_321
timestamp 1666464484
transform 1 0 37296 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_385
timestamp 1666464484
transform 1 0 44464 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_389
timestamp 1666464484
transform 1 0 44912 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_392
timestamp 1666464484
transform 1 0 45248 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_456
timestamp 1666464484
transform 1 0 52416 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_460
timestamp 1666464484
transform 1 0 52864 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_463
timestamp 1666464484
transform 1 0 53200 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_527
timestamp 1666464484
transform 1 0 60368 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_531
timestamp 1666464484
transform 1 0 60816 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_534
timestamp 1666464484
transform 1 0 61152 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_598
timestamp 1666464484
transform 1 0 68320 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_602
timestamp 1666464484
transform 1 0 68768 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_605
timestamp 1666464484
transform 1 0 69104 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_669
timestamp 1666464484
transform 1 0 76272 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_673
timestamp 1666464484
transform 1 0 76720 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_676
timestamp 1666464484
transform 1 0 77056 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_740
timestamp 1666464484
transform 1 0 84224 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_744
timestamp 1666464484
transform 1 0 84672 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_747
timestamp 1666464484
transform 1 0 85008 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_811
timestamp 1666464484
transform 1 0 92176 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_815
timestamp 1666464484
transform 1 0 92624 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_818
timestamp 1666464484
transform 1 0 92960 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_882
timestamp 1666464484
transform 1 0 100128 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_886
timestamp 1666464484
transform 1 0 100576 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_889
timestamp 1666464484
transform 1 0 100912 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_953
timestamp 1666464484
transform 1 0 108080 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_957
timestamp 1666464484
transform 1 0 108528 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_960
timestamp 1666464484
transform 1 0 108864 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1024
timestamp 1666464484
transform 1 0 116032 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1028
timestamp 1666464484
transform 1 0 116480 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_1031
timestamp 1666464484
transform 1 0 116816 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1095
timestamp 1666464484
transform 1 0 123984 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1099
timestamp 1666464484
transform 1 0 124432 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_1102
timestamp 1666464484
transform 1 0 124768 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1166
timestamp 1666464484
transform 1 0 131936 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1170
timestamp 1666464484
transform 1 0 132384 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_1173
timestamp 1666464484
transform 1 0 132720 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1237
timestamp 1666464484
transform 1 0 139888 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1241
timestamp 1666464484
transform 1 0 140336 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_1244
timestamp 1666464484
transform 1 0 140672 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1308
timestamp 1666464484
transform 1 0 147840 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1312
timestamp 1666464484
transform 1 0 148288 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_1315
timestamp 1666464484
transform 1 0 148624 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1379
timestamp 1666464484
transform 1 0 155792 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1383
timestamp 1666464484
transform 1 0 156240 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_1386
timestamp 1666464484
transform 1 0 156576 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1450
timestamp 1666464484
transform 1 0 163744 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1454
timestamp 1666464484
transform 1 0 164192 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_1457
timestamp 1666464484
transform 1 0 164528 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1521
timestamp 1666464484
transform 1 0 171696 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1525
timestamp 1666464484
transform 1 0 172144 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_116_1528
timestamp 1666464484
transform 1 0 172480 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_116_1560
timestamp 1666464484
transform 1 0 176064 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1576
timestamp 1666464484
transform 1 0 177856 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1580
timestamp 1666464484
transform 1 0 178304 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_2
timestamp 1666464484
transform 1 0 1568 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_66
timestamp 1666464484
transform 1 0 8736 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_70
timestamp 1666464484
transform 1 0 9184 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_73
timestamp 1666464484
transform 1 0 9520 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_137
timestamp 1666464484
transform 1 0 16688 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_141
timestamp 1666464484
transform 1 0 17136 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_144
timestamp 1666464484
transform 1 0 17472 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_208
timestamp 1666464484
transform 1 0 24640 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_212
timestamp 1666464484
transform 1 0 25088 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_215
timestamp 1666464484
transform 1 0 25424 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_279
timestamp 1666464484
transform 1 0 32592 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_283
timestamp 1666464484
transform 1 0 33040 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_286
timestamp 1666464484
transform 1 0 33376 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_350
timestamp 1666464484
transform 1 0 40544 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_354
timestamp 1666464484
transform 1 0 40992 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_357
timestamp 1666464484
transform 1 0 41328 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_421
timestamp 1666464484
transform 1 0 48496 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_425
timestamp 1666464484
transform 1 0 48944 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_428
timestamp 1666464484
transform 1 0 49280 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_492
timestamp 1666464484
transform 1 0 56448 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_496
timestamp 1666464484
transform 1 0 56896 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_499
timestamp 1666464484
transform 1 0 57232 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_563
timestamp 1666464484
transform 1 0 64400 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_567
timestamp 1666464484
transform 1 0 64848 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_570
timestamp 1666464484
transform 1 0 65184 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_634
timestamp 1666464484
transform 1 0 72352 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_638
timestamp 1666464484
transform 1 0 72800 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_641
timestamp 1666464484
transform 1 0 73136 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_705
timestamp 1666464484
transform 1 0 80304 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_709
timestamp 1666464484
transform 1 0 80752 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_712
timestamp 1666464484
transform 1 0 81088 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_776
timestamp 1666464484
transform 1 0 88256 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_780
timestamp 1666464484
transform 1 0 88704 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_783
timestamp 1666464484
transform 1 0 89040 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_847
timestamp 1666464484
transform 1 0 96208 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_851
timestamp 1666464484
transform 1 0 96656 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_854
timestamp 1666464484
transform 1 0 96992 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_918
timestamp 1666464484
transform 1 0 104160 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_922
timestamp 1666464484
transform 1 0 104608 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_925
timestamp 1666464484
transform 1 0 104944 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_989
timestamp 1666464484
transform 1 0 112112 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_993
timestamp 1666464484
transform 1 0 112560 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_996
timestamp 1666464484
transform 1 0 112896 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1060
timestamp 1666464484
transform 1 0 120064 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1064
timestamp 1666464484
transform 1 0 120512 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_1067
timestamp 1666464484
transform 1 0 120848 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1131
timestamp 1666464484
transform 1 0 128016 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1135
timestamp 1666464484
transform 1 0 128464 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_1138
timestamp 1666464484
transform 1 0 128800 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1202
timestamp 1666464484
transform 1 0 135968 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1206
timestamp 1666464484
transform 1 0 136416 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_1209
timestamp 1666464484
transform 1 0 136752 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1273
timestamp 1666464484
transform 1 0 143920 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1277
timestamp 1666464484
transform 1 0 144368 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_1280
timestamp 1666464484
transform 1 0 144704 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1344
timestamp 1666464484
transform 1 0 151872 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1348
timestamp 1666464484
transform 1 0 152320 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_1351
timestamp 1666464484
transform 1 0 152656 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1415
timestamp 1666464484
transform 1 0 159824 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1419
timestamp 1666464484
transform 1 0 160272 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_1422
timestamp 1666464484
transform 1 0 160608 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1486
timestamp 1666464484
transform 1 0 167776 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1490
timestamp 1666464484
transform 1 0 168224 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_1493
timestamp 1666464484
transform 1 0 168560 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_1557
timestamp 1666464484
transform 1 0 175728 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1561
timestamp 1666464484
transform 1 0 176176 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_117_1564
timestamp 1666464484
transform 1 0 176512 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1580
timestamp 1666464484
transform 1 0 178304 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_2
timestamp 1666464484
transform 1 0 1568 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_34
timestamp 1666464484
transform 1 0 5152 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_37
timestamp 1666464484
transform 1 0 5488 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_101
timestamp 1666464484
transform 1 0 12656 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_105
timestamp 1666464484
transform 1 0 13104 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_108
timestamp 1666464484
transform 1 0 13440 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_172
timestamp 1666464484
transform 1 0 20608 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_176
timestamp 1666464484
transform 1 0 21056 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_179
timestamp 1666464484
transform 1 0 21392 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_243
timestamp 1666464484
transform 1 0 28560 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_247
timestamp 1666464484
transform 1 0 29008 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_250
timestamp 1666464484
transform 1 0 29344 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_314
timestamp 1666464484
transform 1 0 36512 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_318
timestamp 1666464484
transform 1 0 36960 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_321
timestamp 1666464484
transform 1 0 37296 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_385
timestamp 1666464484
transform 1 0 44464 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_389
timestamp 1666464484
transform 1 0 44912 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_392
timestamp 1666464484
transform 1 0 45248 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_456
timestamp 1666464484
transform 1 0 52416 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_460
timestamp 1666464484
transform 1 0 52864 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_463
timestamp 1666464484
transform 1 0 53200 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_527
timestamp 1666464484
transform 1 0 60368 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_531
timestamp 1666464484
transform 1 0 60816 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_534
timestamp 1666464484
transform 1 0 61152 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_598
timestamp 1666464484
transform 1 0 68320 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_602
timestamp 1666464484
transform 1 0 68768 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_605
timestamp 1666464484
transform 1 0 69104 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_669
timestamp 1666464484
transform 1 0 76272 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_673
timestamp 1666464484
transform 1 0 76720 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_676
timestamp 1666464484
transform 1 0 77056 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_740
timestamp 1666464484
transform 1 0 84224 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_744
timestamp 1666464484
transform 1 0 84672 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_747
timestamp 1666464484
transform 1 0 85008 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_811
timestamp 1666464484
transform 1 0 92176 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_815
timestamp 1666464484
transform 1 0 92624 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_818
timestamp 1666464484
transform 1 0 92960 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_882
timestamp 1666464484
transform 1 0 100128 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_886
timestamp 1666464484
transform 1 0 100576 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_889
timestamp 1666464484
transform 1 0 100912 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_953
timestamp 1666464484
transform 1 0 108080 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_957
timestamp 1666464484
transform 1 0 108528 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_960
timestamp 1666464484
transform 1 0 108864 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1024
timestamp 1666464484
transform 1 0 116032 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1028
timestamp 1666464484
transform 1 0 116480 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_1031
timestamp 1666464484
transform 1 0 116816 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1095
timestamp 1666464484
transform 1 0 123984 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1099
timestamp 1666464484
transform 1 0 124432 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_1102
timestamp 1666464484
transform 1 0 124768 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1166
timestamp 1666464484
transform 1 0 131936 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1170
timestamp 1666464484
transform 1 0 132384 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_1173
timestamp 1666464484
transform 1 0 132720 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1237
timestamp 1666464484
transform 1 0 139888 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1241
timestamp 1666464484
transform 1 0 140336 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_1244
timestamp 1666464484
transform 1 0 140672 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1308
timestamp 1666464484
transform 1 0 147840 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1312
timestamp 1666464484
transform 1 0 148288 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_1315
timestamp 1666464484
transform 1 0 148624 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1379
timestamp 1666464484
transform 1 0 155792 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1383
timestamp 1666464484
transform 1 0 156240 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_1386
timestamp 1666464484
transform 1 0 156576 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1450
timestamp 1666464484
transform 1 0 163744 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1454
timestamp 1666464484
transform 1 0 164192 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_1457
timestamp 1666464484
transform 1 0 164528 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1521
timestamp 1666464484
transform 1 0 171696 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1525
timestamp 1666464484
transform 1 0 172144 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_1528
timestamp 1666464484
transform 1 0 172480 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_118_1560
timestamp 1666464484
transform 1 0 176064 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1576
timestamp 1666464484
transform 1 0 177856 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1580
timestamp 1666464484
transform 1 0 178304 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_2
timestamp 1666464484
transform 1 0 1568 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_66
timestamp 1666464484
transform 1 0 8736 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_70
timestamp 1666464484
transform 1 0 9184 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_73
timestamp 1666464484
transform 1 0 9520 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_137
timestamp 1666464484
transform 1 0 16688 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_141
timestamp 1666464484
transform 1 0 17136 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_144
timestamp 1666464484
transform 1 0 17472 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_208
timestamp 1666464484
transform 1 0 24640 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_212
timestamp 1666464484
transform 1 0 25088 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_215
timestamp 1666464484
transform 1 0 25424 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_279
timestamp 1666464484
transform 1 0 32592 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_283
timestamp 1666464484
transform 1 0 33040 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_286
timestamp 1666464484
transform 1 0 33376 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_350
timestamp 1666464484
transform 1 0 40544 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_354
timestamp 1666464484
transform 1 0 40992 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_357
timestamp 1666464484
transform 1 0 41328 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_421
timestamp 1666464484
transform 1 0 48496 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_425
timestamp 1666464484
transform 1 0 48944 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_428
timestamp 1666464484
transform 1 0 49280 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_492
timestamp 1666464484
transform 1 0 56448 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_496
timestamp 1666464484
transform 1 0 56896 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_499
timestamp 1666464484
transform 1 0 57232 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_563
timestamp 1666464484
transform 1 0 64400 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_567
timestamp 1666464484
transform 1 0 64848 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_570
timestamp 1666464484
transform 1 0 65184 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_634
timestamp 1666464484
transform 1 0 72352 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_638
timestamp 1666464484
transform 1 0 72800 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_641
timestamp 1666464484
transform 1 0 73136 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_705
timestamp 1666464484
transform 1 0 80304 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_709
timestamp 1666464484
transform 1 0 80752 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_712
timestamp 1666464484
transform 1 0 81088 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_776
timestamp 1666464484
transform 1 0 88256 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_780
timestamp 1666464484
transform 1 0 88704 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_783
timestamp 1666464484
transform 1 0 89040 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_847
timestamp 1666464484
transform 1 0 96208 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_851
timestamp 1666464484
transform 1 0 96656 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_854
timestamp 1666464484
transform 1 0 96992 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_918
timestamp 1666464484
transform 1 0 104160 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_922
timestamp 1666464484
transform 1 0 104608 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_925
timestamp 1666464484
transform 1 0 104944 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_989
timestamp 1666464484
transform 1 0 112112 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_993
timestamp 1666464484
transform 1 0 112560 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_996
timestamp 1666464484
transform 1 0 112896 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1060
timestamp 1666464484
transform 1 0 120064 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1064
timestamp 1666464484
transform 1 0 120512 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_1067
timestamp 1666464484
transform 1 0 120848 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1131
timestamp 1666464484
transform 1 0 128016 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1135
timestamp 1666464484
transform 1 0 128464 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_1138
timestamp 1666464484
transform 1 0 128800 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1202
timestamp 1666464484
transform 1 0 135968 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1206
timestamp 1666464484
transform 1 0 136416 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_1209
timestamp 1666464484
transform 1 0 136752 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1273
timestamp 1666464484
transform 1 0 143920 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1277
timestamp 1666464484
transform 1 0 144368 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_1280
timestamp 1666464484
transform 1 0 144704 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1344
timestamp 1666464484
transform 1 0 151872 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1348
timestamp 1666464484
transform 1 0 152320 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_1351
timestamp 1666464484
transform 1 0 152656 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1415
timestamp 1666464484
transform 1 0 159824 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1419
timestamp 1666464484
transform 1 0 160272 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_1422
timestamp 1666464484
transform 1 0 160608 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1486
timestamp 1666464484
transform 1 0 167776 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1490
timestamp 1666464484
transform 1 0 168224 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_1493
timestamp 1666464484
transform 1 0 168560 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_1557
timestamp 1666464484
transform 1 0 175728 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1561
timestamp 1666464484
transform 1 0 176176 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_119_1564
timestamp 1666464484
transform 1 0 176512 0 -1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1580
timestamp 1666464484
transform 1 0 178304 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_120_2
timestamp 1666464484
transform 1 0 1568 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_34
timestamp 1666464484
transform 1 0 5152 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_37
timestamp 1666464484
transform 1 0 5488 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_101
timestamp 1666464484
transform 1 0 12656 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_105
timestamp 1666464484
transform 1 0 13104 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_108
timestamp 1666464484
transform 1 0 13440 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_172
timestamp 1666464484
transform 1 0 20608 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_176
timestamp 1666464484
transform 1 0 21056 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_179
timestamp 1666464484
transform 1 0 21392 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_243
timestamp 1666464484
transform 1 0 28560 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_247
timestamp 1666464484
transform 1 0 29008 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_250
timestamp 1666464484
transform 1 0 29344 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_314
timestamp 1666464484
transform 1 0 36512 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_318
timestamp 1666464484
transform 1 0 36960 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_321
timestamp 1666464484
transform 1 0 37296 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_385
timestamp 1666464484
transform 1 0 44464 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_389
timestamp 1666464484
transform 1 0 44912 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_392
timestamp 1666464484
transform 1 0 45248 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_456
timestamp 1666464484
transform 1 0 52416 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_460
timestamp 1666464484
transform 1 0 52864 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_463
timestamp 1666464484
transform 1 0 53200 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_527
timestamp 1666464484
transform 1 0 60368 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_531
timestamp 1666464484
transform 1 0 60816 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_534
timestamp 1666464484
transform 1 0 61152 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_598
timestamp 1666464484
transform 1 0 68320 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_602
timestamp 1666464484
transform 1 0 68768 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_605
timestamp 1666464484
transform 1 0 69104 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_669
timestamp 1666464484
transform 1 0 76272 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_673
timestamp 1666464484
transform 1 0 76720 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_676
timestamp 1666464484
transform 1 0 77056 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_740
timestamp 1666464484
transform 1 0 84224 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_744
timestamp 1666464484
transform 1 0 84672 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_747
timestamp 1666464484
transform 1 0 85008 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_811
timestamp 1666464484
transform 1 0 92176 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_815
timestamp 1666464484
transform 1 0 92624 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_818
timestamp 1666464484
transform 1 0 92960 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_882
timestamp 1666464484
transform 1 0 100128 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_886
timestamp 1666464484
transform 1 0 100576 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_889
timestamp 1666464484
transform 1 0 100912 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_953
timestamp 1666464484
transform 1 0 108080 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_957
timestamp 1666464484
transform 1 0 108528 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_960
timestamp 1666464484
transform 1 0 108864 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1024
timestamp 1666464484
transform 1 0 116032 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1028
timestamp 1666464484
transform 1 0 116480 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_1031
timestamp 1666464484
transform 1 0 116816 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1095
timestamp 1666464484
transform 1 0 123984 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1099
timestamp 1666464484
transform 1 0 124432 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_1102
timestamp 1666464484
transform 1 0 124768 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1166
timestamp 1666464484
transform 1 0 131936 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1170
timestamp 1666464484
transform 1 0 132384 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_1173
timestamp 1666464484
transform 1 0 132720 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1237
timestamp 1666464484
transform 1 0 139888 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1241
timestamp 1666464484
transform 1 0 140336 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_1244
timestamp 1666464484
transform 1 0 140672 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1308
timestamp 1666464484
transform 1 0 147840 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1312
timestamp 1666464484
transform 1 0 148288 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_1315
timestamp 1666464484
transform 1 0 148624 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1379
timestamp 1666464484
transform 1 0 155792 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1383
timestamp 1666464484
transform 1 0 156240 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_1386
timestamp 1666464484
transform 1 0 156576 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1450
timestamp 1666464484
transform 1 0 163744 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1454
timestamp 1666464484
transform 1 0 164192 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_1457
timestamp 1666464484
transform 1 0 164528 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1521
timestamp 1666464484
transform 1 0 171696 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1525
timestamp 1666464484
transform 1 0 172144 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_120_1528
timestamp 1666464484
transform 1 0 172480 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_120_1560
timestamp 1666464484
transform 1 0 176064 0 1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1576
timestamp 1666464484
transform 1 0 177856 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1580
timestamp 1666464484
transform 1 0 178304 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_2
timestamp 1666464484
transform 1 0 1568 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_66
timestamp 1666464484
transform 1 0 8736 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_70
timestamp 1666464484
transform 1 0 9184 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_73
timestamp 1666464484
transform 1 0 9520 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_137
timestamp 1666464484
transform 1 0 16688 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_141
timestamp 1666464484
transform 1 0 17136 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_144
timestamp 1666464484
transform 1 0 17472 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_208
timestamp 1666464484
transform 1 0 24640 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_212
timestamp 1666464484
transform 1 0 25088 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_215
timestamp 1666464484
transform 1 0 25424 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_279
timestamp 1666464484
transform 1 0 32592 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_283
timestamp 1666464484
transform 1 0 33040 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_286
timestamp 1666464484
transform 1 0 33376 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_350
timestamp 1666464484
transform 1 0 40544 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_354
timestamp 1666464484
transform 1 0 40992 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_357
timestamp 1666464484
transform 1 0 41328 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_421
timestamp 1666464484
transform 1 0 48496 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_425
timestamp 1666464484
transform 1 0 48944 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_428
timestamp 1666464484
transform 1 0 49280 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_492
timestamp 1666464484
transform 1 0 56448 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_496
timestamp 1666464484
transform 1 0 56896 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_499
timestamp 1666464484
transform 1 0 57232 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_563
timestamp 1666464484
transform 1 0 64400 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_567
timestamp 1666464484
transform 1 0 64848 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_570
timestamp 1666464484
transform 1 0 65184 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_634
timestamp 1666464484
transform 1 0 72352 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_638
timestamp 1666464484
transform 1 0 72800 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_641
timestamp 1666464484
transform 1 0 73136 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_705
timestamp 1666464484
transform 1 0 80304 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_709
timestamp 1666464484
transform 1 0 80752 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_712
timestamp 1666464484
transform 1 0 81088 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_776
timestamp 1666464484
transform 1 0 88256 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_780
timestamp 1666464484
transform 1 0 88704 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_783
timestamp 1666464484
transform 1 0 89040 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_847
timestamp 1666464484
transform 1 0 96208 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_851
timestamp 1666464484
transform 1 0 96656 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_854
timestamp 1666464484
transform 1 0 96992 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_918
timestamp 1666464484
transform 1 0 104160 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_922
timestamp 1666464484
transform 1 0 104608 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_925
timestamp 1666464484
transform 1 0 104944 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_989
timestamp 1666464484
transform 1 0 112112 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_993
timestamp 1666464484
transform 1 0 112560 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_996
timestamp 1666464484
transform 1 0 112896 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1060
timestamp 1666464484
transform 1 0 120064 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1064
timestamp 1666464484
transform 1 0 120512 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_1067
timestamp 1666464484
transform 1 0 120848 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1131
timestamp 1666464484
transform 1 0 128016 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1135
timestamp 1666464484
transform 1 0 128464 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_1138
timestamp 1666464484
transform 1 0 128800 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1202
timestamp 1666464484
transform 1 0 135968 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1206
timestamp 1666464484
transform 1 0 136416 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_1209
timestamp 1666464484
transform 1 0 136752 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1273
timestamp 1666464484
transform 1 0 143920 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1277
timestamp 1666464484
transform 1 0 144368 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_1280
timestamp 1666464484
transform 1 0 144704 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1344
timestamp 1666464484
transform 1 0 151872 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1348
timestamp 1666464484
transform 1 0 152320 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_1351
timestamp 1666464484
transform 1 0 152656 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1415
timestamp 1666464484
transform 1 0 159824 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1419
timestamp 1666464484
transform 1 0 160272 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_1422
timestamp 1666464484
transform 1 0 160608 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1486
timestamp 1666464484
transform 1 0 167776 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1490
timestamp 1666464484
transform 1 0 168224 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_1493
timestamp 1666464484
transform 1 0 168560 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1557
timestamp 1666464484
transform 1 0 175728 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1561
timestamp 1666464484
transform 1 0 176176 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_121_1564
timestamp 1666464484
transform 1 0 176512 0 -1 98784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1580
timestamp 1666464484
transform 1 0 178304 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_122_2
timestamp 1666464484
transform 1 0 1568 0 1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_34
timestamp 1666464484
transform 1 0 5152 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_37
timestamp 1666464484
transform 1 0 5488 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_101
timestamp 1666464484
transform 1 0 12656 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_105
timestamp 1666464484
transform 1 0 13104 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_108
timestamp 1666464484
transform 1 0 13440 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_172
timestamp 1666464484
transform 1 0 20608 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_176
timestamp 1666464484
transform 1 0 21056 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_179
timestamp 1666464484
transform 1 0 21392 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_243
timestamp 1666464484
transform 1 0 28560 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_247
timestamp 1666464484
transform 1 0 29008 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_250
timestamp 1666464484
transform 1 0 29344 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_314
timestamp 1666464484
transform 1 0 36512 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_318
timestamp 1666464484
transform 1 0 36960 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_321
timestamp 1666464484
transform 1 0 37296 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_385
timestamp 1666464484
transform 1 0 44464 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_389
timestamp 1666464484
transform 1 0 44912 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_392
timestamp 1666464484
transform 1 0 45248 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_456
timestamp 1666464484
transform 1 0 52416 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_460
timestamp 1666464484
transform 1 0 52864 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_463
timestamp 1666464484
transform 1 0 53200 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_527
timestamp 1666464484
transform 1 0 60368 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_531
timestamp 1666464484
transform 1 0 60816 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_534
timestamp 1666464484
transform 1 0 61152 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_598
timestamp 1666464484
transform 1 0 68320 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_602
timestamp 1666464484
transform 1 0 68768 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_605
timestamp 1666464484
transform 1 0 69104 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_669
timestamp 1666464484
transform 1 0 76272 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_673
timestamp 1666464484
transform 1 0 76720 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_676
timestamp 1666464484
transform 1 0 77056 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_740
timestamp 1666464484
transform 1 0 84224 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_744
timestamp 1666464484
transform 1 0 84672 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_747
timestamp 1666464484
transform 1 0 85008 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_811
timestamp 1666464484
transform 1 0 92176 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_815
timestamp 1666464484
transform 1 0 92624 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_818
timestamp 1666464484
transform 1 0 92960 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_882
timestamp 1666464484
transform 1 0 100128 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_886
timestamp 1666464484
transform 1 0 100576 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_889
timestamp 1666464484
transform 1 0 100912 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_953
timestamp 1666464484
transform 1 0 108080 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_957
timestamp 1666464484
transform 1 0 108528 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_960
timestamp 1666464484
transform 1 0 108864 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1024
timestamp 1666464484
transform 1 0 116032 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1028
timestamp 1666464484
transform 1 0 116480 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_1031
timestamp 1666464484
transform 1 0 116816 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1095
timestamp 1666464484
transform 1 0 123984 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1099
timestamp 1666464484
transform 1 0 124432 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_1102
timestamp 1666464484
transform 1 0 124768 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1166
timestamp 1666464484
transform 1 0 131936 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1170
timestamp 1666464484
transform 1 0 132384 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_1173
timestamp 1666464484
transform 1 0 132720 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1237
timestamp 1666464484
transform 1 0 139888 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1241
timestamp 1666464484
transform 1 0 140336 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_1244
timestamp 1666464484
transform 1 0 140672 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1308
timestamp 1666464484
transform 1 0 147840 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1312
timestamp 1666464484
transform 1 0 148288 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_1315
timestamp 1666464484
transform 1 0 148624 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1379
timestamp 1666464484
transform 1 0 155792 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1383
timestamp 1666464484
transform 1 0 156240 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_1386
timestamp 1666464484
transform 1 0 156576 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1450
timestamp 1666464484
transform 1 0 163744 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1454
timestamp 1666464484
transform 1 0 164192 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_1457
timestamp 1666464484
transform 1 0 164528 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1521
timestamp 1666464484
transform 1 0 171696 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1525
timestamp 1666464484
transform 1 0 172144 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_122_1528
timestamp 1666464484
transform 1 0 172480 0 1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_122_1560
timestamp 1666464484
transform 1 0 176064 0 1 98784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1576
timestamp 1666464484
transform 1 0 177856 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1580
timestamp 1666464484
transform 1 0 178304 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_2
timestamp 1666464484
transform 1 0 1568 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_66
timestamp 1666464484
transform 1 0 8736 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_70
timestamp 1666464484
transform 1 0 9184 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_73
timestamp 1666464484
transform 1 0 9520 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_137
timestamp 1666464484
transform 1 0 16688 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_141
timestamp 1666464484
transform 1 0 17136 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_144
timestamp 1666464484
transform 1 0 17472 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_208
timestamp 1666464484
transform 1 0 24640 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_212
timestamp 1666464484
transform 1 0 25088 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_215
timestamp 1666464484
transform 1 0 25424 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_279
timestamp 1666464484
transform 1 0 32592 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_283
timestamp 1666464484
transform 1 0 33040 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_286
timestamp 1666464484
transform 1 0 33376 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_350
timestamp 1666464484
transform 1 0 40544 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_354
timestamp 1666464484
transform 1 0 40992 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_357
timestamp 1666464484
transform 1 0 41328 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_421
timestamp 1666464484
transform 1 0 48496 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_425
timestamp 1666464484
transform 1 0 48944 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_428
timestamp 1666464484
transform 1 0 49280 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_492
timestamp 1666464484
transform 1 0 56448 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_496
timestamp 1666464484
transform 1 0 56896 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_499
timestamp 1666464484
transform 1 0 57232 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_563
timestamp 1666464484
transform 1 0 64400 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_567
timestamp 1666464484
transform 1 0 64848 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_570
timestamp 1666464484
transform 1 0 65184 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_634
timestamp 1666464484
transform 1 0 72352 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_638
timestamp 1666464484
transform 1 0 72800 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_641
timestamp 1666464484
transform 1 0 73136 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_705
timestamp 1666464484
transform 1 0 80304 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_709
timestamp 1666464484
transform 1 0 80752 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_712
timestamp 1666464484
transform 1 0 81088 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_776
timestamp 1666464484
transform 1 0 88256 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_780
timestamp 1666464484
transform 1 0 88704 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_783
timestamp 1666464484
transform 1 0 89040 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_847
timestamp 1666464484
transform 1 0 96208 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_851
timestamp 1666464484
transform 1 0 96656 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_854
timestamp 1666464484
transform 1 0 96992 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_918
timestamp 1666464484
transform 1 0 104160 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_922
timestamp 1666464484
transform 1 0 104608 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_925
timestamp 1666464484
transform 1 0 104944 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_989
timestamp 1666464484
transform 1 0 112112 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_993
timestamp 1666464484
transform 1 0 112560 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_996
timestamp 1666464484
transform 1 0 112896 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1060
timestamp 1666464484
transform 1 0 120064 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1064
timestamp 1666464484
transform 1 0 120512 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_1067
timestamp 1666464484
transform 1 0 120848 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1131
timestamp 1666464484
transform 1 0 128016 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1135
timestamp 1666464484
transform 1 0 128464 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_1138
timestamp 1666464484
transform 1 0 128800 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1202
timestamp 1666464484
transform 1 0 135968 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1206
timestamp 1666464484
transform 1 0 136416 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_1209
timestamp 1666464484
transform 1 0 136752 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1273
timestamp 1666464484
transform 1 0 143920 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1277
timestamp 1666464484
transform 1 0 144368 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_1280
timestamp 1666464484
transform 1 0 144704 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1344
timestamp 1666464484
transform 1 0 151872 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1348
timestamp 1666464484
transform 1 0 152320 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_1351
timestamp 1666464484
transform 1 0 152656 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1415
timestamp 1666464484
transform 1 0 159824 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1419
timestamp 1666464484
transform 1 0 160272 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_1422
timestamp 1666464484
transform 1 0 160608 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1486
timestamp 1666464484
transform 1 0 167776 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1490
timestamp 1666464484
transform 1 0 168224 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_1493
timestamp 1666464484
transform 1 0 168560 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_1557
timestamp 1666464484
transform 1 0 175728 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1561
timestamp 1666464484
transform 1 0 176176 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_123_1564
timestamp 1666464484
transform 1 0 176512 0 -1 100352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1580
timestamp 1666464484
transform 1 0 178304 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_124_2
timestamp 1666464484
transform 1 0 1568 0 1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_34
timestamp 1666464484
transform 1 0 5152 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_37
timestamp 1666464484
transform 1 0 5488 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_101
timestamp 1666464484
transform 1 0 12656 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_105
timestamp 1666464484
transform 1 0 13104 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_108
timestamp 1666464484
transform 1 0 13440 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_172
timestamp 1666464484
transform 1 0 20608 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_176
timestamp 1666464484
transform 1 0 21056 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_179
timestamp 1666464484
transform 1 0 21392 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_243
timestamp 1666464484
transform 1 0 28560 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_247
timestamp 1666464484
transform 1 0 29008 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_250
timestamp 1666464484
transform 1 0 29344 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_314
timestamp 1666464484
transform 1 0 36512 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_318
timestamp 1666464484
transform 1 0 36960 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_321
timestamp 1666464484
transform 1 0 37296 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_385
timestamp 1666464484
transform 1 0 44464 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_389
timestamp 1666464484
transform 1 0 44912 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_392
timestamp 1666464484
transform 1 0 45248 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_456
timestamp 1666464484
transform 1 0 52416 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_460
timestamp 1666464484
transform 1 0 52864 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_463
timestamp 1666464484
transform 1 0 53200 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_527
timestamp 1666464484
transform 1 0 60368 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_531
timestamp 1666464484
transform 1 0 60816 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_534
timestamp 1666464484
transform 1 0 61152 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_598
timestamp 1666464484
transform 1 0 68320 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_602
timestamp 1666464484
transform 1 0 68768 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_605
timestamp 1666464484
transform 1 0 69104 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_669
timestamp 1666464484
transform 1 0 76272 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_673
timestamp 1666464484
transform 1 0 76720 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_676
timestamp 1666464484
transform 1 0 77056 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_740
timestamp 1666464484
transform 1 0 84224 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_744
timestamp 1666464484
transform 1 0 84672 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_747
timestamp 1666464484
transform 1 0 85008 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_811
timestamp 1666464484
transform 1 0 92176 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_815
timestamp 1666464484
transform 1 0 92624 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_818
timestamp 1666464484
transform 1 0 92960 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_882
timestamp 1666464484
transform 1 0 100128 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_886
timestamp 1666464484
transform 1 0 100576 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_889
timestamp 1666464484
transform 1 0 100912 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_953
timestamp 1666464484
transform 1 0 108080 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_957
timestamp 1666464484
transform 1 0 108528 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_960
timestamp 1666464484
transform 1 0 108864 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1024
timestamp 1666464484
transform 1 0 116032 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1028
timestamp 1666464484
transform 1 0 116480 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_1031
timestamp 1666464484
transform 1 0 116816 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1095
timestamp 1666464484
transform 1 0 123984 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1099
timestamp 1666464484
transform 1 0 124432 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_1102
timestamp 1666464484
transform 1 0 124768 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1166
timestamp 1666464484
transform 1 0 131936 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1170
timestamp 1666464484
transform 1 0 132384 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_1173
timestamp 1666464484
transform 1 0 132720 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1237
timestamp 1666464484
transform 1 0 139888 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1241
timestamp 1666464484
transform 1 0 140336 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_1244
timestamp 1666464484
transform 1 0 140672 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1308
timestamp 1666464484
transform 1 0 147840 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1312
timestamp 1666464484
transform 1 0 148288 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_1315
timestamp 1666464484
transform 1 0 148624 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1379
timestamp 1666464484
transform 1 0 155792 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1383
timestamp 1666464484
transform 1 0 156240 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_1386
timestamp 1666464484
transform 1 0 156576 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1450
timestamp 1666464484
transform 1 0 163744 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1454
timestamp 1666464484
transform 1 0 164192 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_1457
timestamp 1666464484
transform 1 0 164528 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1521
timestamp 1666464484
transform 1 0 171696 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1525
timestamp 1666464484
transform 1 0 172144 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_124_1528
timestamp 1666464484
transform 1 0 172480 0 1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_124_1560
timestamp 1666464484
transform 1 0 176064 0 1 100352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1576
timestamp 1666464484
transform 1 0 177856 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1580
timestamp 1666464484
transform 1 0 178304 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_2
timestamp 1666464484
transform 1 0 1568 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_66
timestamp 1666464484
transform 1 0 8736 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_70
timestamp 1666464484
transform 1 0 9184 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_73
timestamp 1666464484
transform 1 0 9520 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_137
timestamp 1666464484
transform 1 0 16688 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_141
timestamp 1666464484
transform 1 0 17136 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_144
timestamp 1666464484
transform 1 0 17472 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_208
timestamp 1666464484
transform 1 0 24640 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_212
timestamp 1666464484
transform 1 0 25088 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_215
timestamp 1666464484
transform 1 0 25424 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_279
timestamp 1666464484
transform 1 0 32592 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_283
timestamp 1666464484
transform 1 0 33040 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_286
timestamp 1666464484
transform 1 0 33376 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_350
timestamp 1666464484
transform 1 0 40544 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_354
timestamp 1666464484
transform 1 0 40992 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_357
timestamp 1666464484
transform 1 0 41328 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_421
timestamp 1666464484
transform 1 0 48496 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_425
timestamp 1666464484
transform 1 0 48944 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_428
timestamp 1666464484
transform 1 0 49280 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_492
timestamp 1666464484
transform 1 0 56448 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_496
timestamp 1666464484
transform 1 0 56896 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_499
timestamp 1666464484
transform 1 0 57232 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_563
timestamp 1666464484
transform 1 0 64400 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_567
timestamp 1666464484
transform 1 0 64848 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_570
timestamp 1666464484
transform 1 0 65184 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_634
timestamp 1666464484
transform 1 0 72352 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_638
timestamp 1666464484
transform 1 0 72800 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_641
timestamp 1666464484
transform 1 0 73136 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_705
timestamp 1666464484
transform 1 0 80304 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_709
timestamp 1666464484
transform 1 0 80752 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_712
timestamp 1666464484
transform 1 0 81088 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_776
timestamp 1666464484
transform 1 0 88256 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_780
timestamp 1666464484
transform 1 0 88704 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_783
timestamp 1666464484
transform 1 0 89040 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_847
timestamp 1666464484
transform 1 0 96208 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_851
timestamp 1666464484
transform 1 0 96656 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_854
timestamp 1666464484
transform 1 0 96992 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_918
timestamp 1666464484
transform 1 0 104160 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_922
timestamp 1666464484
transform 1 0 104608 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_925
timestamp 1666464484
transform 1 0 104944 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_989
timestamp 1666464484
transform 1 0 112112 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_993
timestamp 1666464484
transform 1 0 112560 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_996
timestamp 1666464484
transform 1 0 112896 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1060
timestamp 1666464484
transform 1 0 120064 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1064
timestamp 1666464484
transform 1 0 120512 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_1067
timestamp 1666464484
transform 1 0 120848 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1131
timestamp 1666464484
transform 1 0 128016 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1135
timestamp 1666464484
transform 1 0 128464 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_1138
timestamp 1666464484
transform 1 0 128800 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1202
timestamp 1666464484
transform 1 0 135968 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1206
timestamp 1666464484
transform 1 0 136416 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_1209
timestamp 1666464484
transform 1 0 136752 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1273
timestamp 1666464484
transform 1 0 143920 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1277
timestamp 1666464484
transform 1 0 144368 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_1280
timestamp 1666464484
transform 1 0 144704 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1344
timestamp 1666464484
transform 1 0 151872 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1348
timestamp 1666464484
transform 1 0 152320 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_1351
timestamp 1666464484
transform 1 0 152656 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1415
timestamp 1666464484
transform 1 0 159824 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1419
timestamp 1666464484
transform 1 0 160272 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_1422
timestamp 1666464484
transform 1 0 160608 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1486
timestamp 1666464484
transform 1 0 167776 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1490
timestamp 1666464484
transform 1 0 168224 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_1493
timestamp 1666464484
transform 1 0 168560 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_1557
timestamp 1666464484
transform 1 0 175728 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1561
timestamp 1666464484
transform 1 0 176176 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_125_1564
timestamp 1666464484
transform 1 0 176512 0 -1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1580
timestamp 1666464484
transform 1 0 178304 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_126_2
timestamp 1666464484
transform 1 0 1568 0 1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_34
timestamp 1666464484
transform 1 0 5152 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_37
timestamp 1666464484
transform 1 0 5488 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_101
timestamp 1666464484
transform 1 0 12656 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_105
timestamp 1666464484
transform 1 0 13104 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_108
timestamp 1666464484
transform 1 0 13440 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_172
timestamp 1666464484
transform 1 0 20608 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_176
timestamp 1666464484
transform 1 0 21056 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_179
timestamp 1666464484
transform 1 0 21392 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_243
timestamp 1666464484
transform 1 0 28560 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_247
timestamp 1666464484
transform 1 0 29008 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_250
timestamp 1666464484
transform 1 0 29344 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_314
timestamp 1666464484
transform 1 0 36512 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_318
timestamp 1666464484
transform 1 0 36960 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_321
timestamp 1666464484
transform 1 0 37296 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_385
timestamp 1666464484
transform 1 0 44464 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_389
timestamp 1666464484
transform 1 0 44912 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_392
timestamp 1666464484
transform 1 0 45248 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_456
timestamp 1666464484
transform 1 0 52416 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_460
timestamp 1666464484
transform 1 0 52864 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_463
timestamp 1666464484
transform 1 0 53200 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_527
timestamp 1666464484
transform 1 0 60368 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_531
timestamp 1666464484
transform 1 0 60816 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_534
timestamp 1666464484
transform 1 0 61152 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_598
timestamp 1666464484
transform 1 0 68320 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_602
timestamp 1666464484
transform 1 0 68768 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_605
timestamp 1666464484
transform 1 0 69104 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_669
timestamp 1666464484
transform 1 0 76272 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_673
timestamp 1666464484
transform 1 0 76720 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_676
timestamp 1666464484
transform 1 0 77056 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_740
timestamp 1666464484
transform 1 0 84224 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_744
timestamp 1666464484
transform 1 0 84672 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_747
timestamp 1666464484
transform 1 0 85008 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_811
timestamp 1666464484
transform 1 0 92176 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_815
timestamp 1666464484
transform 1 0 92624 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_818
timestamp 1666464484
transform 1 0 92960 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_882
timestamp 1666464484
transform 1 0 100128 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_886
timestamp 1666464484
transform 1 0 100576 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_889
timestamp 1666464484
transform 1 0 100912 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_953
timestamp 1666464484
transform 1 0 108080 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_957
timestamp 1666464484
transform 1 0 108528 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_960
timestamp 1666464484
transform 1 0 108864 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1024
timestamp 1666464484
transform 1 0 116032 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1028
timestamp 1666464484
transform 1 0 116480 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_1031
timestamp 1666464484
transform 1 0 116816 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1095
timestamp 1666464484
transform 1 0 123984 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1099
timestamp 1666464484
transform 1 0 124432 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_1102
timestamp 1666464484
transform 1 0 124768 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1166
timestamp 1666464484
transform 1 0 131936 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1170
timestamp 1666464484
transform 1 0 132384 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_1173
timestamp 1666464484
transform 1 0 132720 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1237
timestamp 1666464484
transform 1 0 139888 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1241
timestamp 1666464484
transform 1 0 140336 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_1244
timestamp 1666464484
transform 1 0 140672 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1308
timestamp 1666464484
transform 1 0 147840 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1312
timestamp 1666464484
transform 1 0 148288 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_1315
timestamp 1666464484
transform 1 0 148624 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1379
timestamp 1666464484
transform 1 0 155792 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1383
timestamp 1666464484
transform 1 0 156240 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_1386
timestamp 1666464484
transform 1 0 156576 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1450
timestamp 1666464484
transform 1 0 163744 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1454
timestamp 1666464484
transform 1 0 164192 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_1457
timestamp 1666464484
transform 1 0 164528 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1521
timestamp 1666464484
transform 1 0 171696 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1525
timestamp 1666464484
transform 1 0 172144 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_126_1528
timestamp 1666464484
transform 1 0 172480 0 1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_126_1560
timestamp 1666464484
transform 1 0 176064 0 1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1576
timestamp 1666464484
transform 1 0 177856 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1580
timestamp 1666464484
transform 1 0 178304 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_2
timestamp 1666464484
transform 1 0 1568 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_66
timestamp 1666464484
transform 1 0 8736 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_70
timestamp 1666464484
transform 1 0 9184 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_73
timestamp 1666464484
transform 1 0 9520 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_137
timestamp 1666464484
transform 1 0 16688 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_141
timestamp 1666464484
transform 1 0 17136 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_144
timestamp 1666464484
transform 1 0 17472 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_208
timestamp 1666464484
transform 1 0 24640 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_212
timestamp 1666464484
transform 1 0 25088 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_215
timestamp 1666464484
transform 1 0 25424 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_279
timestamp 1666464484
transform 1 0 32592 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_283
timestamp 1666464484
transform 1 0 33040 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_286
timestamp 1666464484
transform 1 0 33376 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_350
timestamp 1666464484
transform 1 0 40544 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_354
timestamp 1666464484
transform 1 0 40992 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_357
timestamp 1666464484
transform 1 0 41328 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_421
timestamp 1666464484
transform 1 0 48496 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_425
timestamp 1666464484
transform 1 0 48944 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_428
timestamp 1666464484
transform 1 0 49280 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_492
timestamp 1666464484
transform 1 0 56448 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_496
timestamp 1666464484
transform 1 0 56896 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_499
timestamp 1666464484
transform 1 0 57232 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_563
timestamp 1666464484
transform 1 0 64400 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_567
timestamp 1666464484
transform 1 0 64848 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_570
timestamp 1666464484
transform 1 0 65184 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_634
timestamp 1666464484
transform 1 0 72352 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_638
timestamp 1666464484
transform 1 0 72800 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_641
timestamp 1666464484
transform 1 0 73136 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_705
timestamp 1666464484
transform 1 0 80304 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_709
timestamp 1666464484
transform 1 0 80752 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_712
timestamp 1666464484
transform 1 0 81088 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_776
timestamp 1666464484
transform 1 0 88256 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_780
timestamp 1666464484
transform 1 0 88704 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_783
timestamp 1666464484
transform 1 0 89040 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_847
timestamp 1666464484
transform 1 0 96208 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_851
timestamp 1666464484
transform 1 0 96656 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_854
timestamp 1666464484
transform 1 0 96992 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_918
timestamp 1666464484
transform 1 0 104160 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_922
timestamp 1666464484
transform 1 0 104608 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_925
timestamp 1666464484
transform 1 0 104944 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_989
timestamp 1666464484
transform 1 0 112112 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_993
timestamp 1666464484
transform 1 0 112560 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_996
timestamp 1666464484
transform 1 0 112896 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1060
timestamp 1666464484
transform 1 0 120064 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1064
timestamp 1666464484
transform 1 0 120512 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_1067
timestamp 1666464484
transform 1 0 120848 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1131
timestamp 1666464484
transform 1 0 128016 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1135
timestamp 1666464484
transform 1 0 128464 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_1138
timestamp 1666464484
transform 1 0 128800 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1202
timestamp 1666464484
transform 1 0 135968 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1206
timestamp 1666464484
transform 1 0 136416 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_1209
timestamp 1666464484
transform 1 0 136752 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1273
timestamp 1666464484
transform 1 0 143920 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1277
timestamp 1666464484
transform 1 0 144368 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_1280
timestamp 1666464484
transform 1 0 144704 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1344
timestamp 1666464484
transform 1 0 151872 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1348
timestamp 1666464484
transform 1 0 152320 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_1351
timestamp 1666464484
transform 1 0 152656 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1415
timestamp 1666464484
transform 1 0 159824 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1419
timestamp 1666464484
transform 1 0 160272 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_1422
timestamp 1666464484
transform 1 0 160608 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1486
timestamp 1666464484
transform 1 0 167776 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1490
timestamp 1666464484
transform 1 0 168224 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_1493
timestamp 1666464484
transform 1 0 168560 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1557
timestamp 1666464484
transform 1 0 175728 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1561
timestamp 1666464484
transform 1 0 176176 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_127_1564
timestamp 1666464484
transform 1 0 176512 0 -1 103488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1580
timestamp 1666464484
transform 1 0 178304 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_128_2
timestamp 1666464484
transform 1 0 1568 0 1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_34
timestamp 1666464484
transform 1 0 5152 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_37
timestamp 1666464484
transform 1 0 5488 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_101
timestamp 1666464484
transform 1 0 12656 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_105
timestamp 1666464484
transform 1 0 13104 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_108
timestamp 1666464484
transform 1 0 13440 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_172
timestamp 1666464484
transform 1 0 20608 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_176
timestamp 1666464484
transform 1 0 21056 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_179
timestamp 1666464484
transform 1 0 21392 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_243
timestamp 1666464484
transform 1 0 28560 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_247
timestamp 1666464484
transform 1 0 29008 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_250
timestamp 1666464484
transform 1 0 29344 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_314
timestamp 1666464484
transform 1 0 36512 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_318
timestamp 1666464484
transform 1 0 36960 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_321
timestamp 1666464484
transform 1 0 37296 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_385
timestamp 1666464484
transform 1 0 44464 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_389
timestamp 1666464484
transform 1 0 44912 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_392
timestamp 1666464484
transform 1 0 45248 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_456
timestamp 1666464484
transform 1 0 52416 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_460
timestamp 1666464484
transform 1 0 52864 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_463
timestamp 1666464484
transform 1 0 53200 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_527
timestamp 1666464484
transform 1 0 60368 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_531
timestamp 1666464484
transform 1 0 60816 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_534
timestamp 1666464484
transform 1 0 61152 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_598
timestamp 1666464484
transform 1 0 68320 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_602
timestamp 1666464484
transform 1 0 68768 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_605
timestamp 1666464484
transform 1 0 69104 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_669
timestamp 1666464484
transform 1 0 76272 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_673
timestamp 1666464484
transform 1 0 76720 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_676
timestamp 1666464484
transform 1 0 77056 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_740
timestamp 1666464484
transform 1 0 84224 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_744
timestamp 1666464484
transform 1 0 84672 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_747
timestamp 1666464484
transform 1 0 85008 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_811
timestamp 1666464484
transform 1 0 92176 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_815
timestamp 1666464484
transform 1 0 92624 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_818
timestamp 1666464484
transform 1 0 92960 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_882
timestamp 1666464484
transform 1 0 100128 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_886
timestamp 1666464484
transform 1 0 100576 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_889
timestamp 1666464484
transform 1 0 100912 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_953
timestamp 1666464484
transform 1 0 108080 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_957
timestamp 1666464484
transform 1 0 108528 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_960
timestamp 1666464484
transform 1 0 108864 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1024
timestamp 1666464484
transform 1 0 116032 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1028
timestamp 1666464484
transform 1 0 116480 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_1031
timestamp 1666464484
transform 1 0 116816 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1095
timestamp 1666464484
transform 1 0 123984 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1099
timestamp 1666464484
transform 1 0 124432 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_1102
timestamp 1666464484
transform 1 0 124768 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1166
timestamp 1666464484
transform 1 0 131936 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1170
timestamp 1666464484
transform 1 0 132384 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_1173
timestamp 1666464484
transform 1 0 132720 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1237
timestamp 1666464484
transform 1 0 139888 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1241
timestamp 1666464484
transform 1 0 140336 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_1244
timestamp 1666464484
transform 1 0 140672 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1308
timestamp 1666464484
transform 1 0 147840 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1312
timestamp 1666464484
transform 1 0 148288 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_1315
timestamp 1666464484
transform 1 0 148624 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1379
timestamp 1666464484
transform 1 0 155792 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1383
timestamp 1666464484
transform 1 0 156240 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_1386
timestamp 1666464484
transform 1 0 156576 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1450
timestamp 1666464484
transform 1 0 163744 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1454
timestamp 1666464484
transform 1 0 164192 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_1457
timestamp 1666464484
transform 1 0 164528 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1521
timestamp 1666464484
transform 1 0 171696 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1525
timestamp 1666464484
transform 1 0 172144 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_128_1528
timestamp 1666464484
transform 1 0 172480 0 1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_128_1560
timestamp 1666464484
transform 1 0 176064 0 1 103488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1576
timestamp 1666464484
transform 1 0 177856 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1580
timestamp 1666464484
transform 1 0 178304 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_2
timestamp 1666464484
transform 1 0 1568 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_66
timestamp 1666464484
transform 1 0 8736 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_70
timestamp 1666464484
transform 1 0 9184 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_73
timestamp 1666464484
transform 1 0 9520 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_137
timestamp 1666464484
transform 1 0 16688 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_141
timestamp 1666464484
transform 1 0 17136 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_144
timestamp 1666464484
transform 1 0 17472 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_208
timestamp 1666464484
transform 1 0 24640 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_212
timestamp 1666464484
transform 1 0 25088 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_215
timestamp 1666464484
transform 1 0 25424 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_279
timestamp 1666464484
transform 1 0 32592 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_283
timestamp 1666464484
transform 1 0 33040 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_286
timestamp 1666464484
transform 1 0 33376 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_350
timestamp 1666464484
transform 1 0 40544 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_354
timestamp 1666464484
transform 1 0 40992 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_357
timestamp 1666464484
transform 1 0 41328 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_421
timestamp 1666464484
transform 1 0 48496 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_425
timestamp 1666464484
transform 1 0 48944 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_428
timestamp 1666464484
transform 1 0 49280 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_492
timestamp 1666464484
transform 1 0 56448 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_496
timestamp 1666464484
transform 1 0 56896 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_499
timestamp 1666464484
transform 1 0 57232 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_563
timestamp 1666464484
transform 1 0 64400 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_567
timestamp 1666464484
transform 1 0 64848 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_570
timestamp 1666464484
transform 1 0 65184 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_634
timestamp 1666464484
transform 1 0 72352 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_638
timestamp 1666464484
transform 1 0 72800 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_641
timestamp 1666464484
transform 1 0 73136 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_705
timestamp 1666464484
transform 1 0 80304 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_709
timestamp 1666464484
transform 1 0 80752 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_712
timestamp 1666464484
transform 1 0 81088 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_776
timestamp 1666464484
transform 1 0 88256 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_780
timestamp 1666464484
transform 1 0 88704 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_783
timestamp 1666464484
transform 1 0 89040 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_847
timestamp 1666464484
transform 1 0 96208 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_851
timestamp 1666464484
transform 1 0 96656 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_854
timestamp 1666464484
transform 1 0 96992 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_918
timestamp 1666464484
transform 1 0 104160 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_922
timestamp 1666464484
transform 1 0 104608 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_925
timestamp 1666464484
transform 1 0 104944 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_989
timestamp 1666464484
transform 1 0 112112 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_993
timestamp 1666464484
transform 1 0 112560 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_996
timestamp 1666464484
transform 1 0 112896 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1060
timestamp 1666464484
transform 1 0 120064 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1064
timestamp 1666464484
transform 1 0 120512 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_1067
timestamp 1666464484
transform 1 0 120848 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1131
timestamp 1666464484
transform 1 0 128016 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1135
timestamp 1666464484
transform 1 0 128464 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_1138
timestamp 1666464484
transform 1 0 128800 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1202
timestamp 1666464484
transform 1 0 135968 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1206
timestamp 1666464484
transform 1 0 136416 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_1209
timestamp 1666464484
transform 1 0 136752 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1273
timestamp 1666464484
transform 1 0 143920 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1277
timestamp 1666464484
transform 1 0 144368 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_1280
timestamp 1666464484
transform 1 0 144704 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1344
timestamp 1666464484
transform 1 0 151872 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1348
timestamp 1666464484
transform 1 0 152320 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_1351
timestamp 1666464484
transform 1 0 152656 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1415
timestamp 1666464484
transform 1 0 159824 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1419
timestamp 1666464484
transform 1 0 160272 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_1422
timestamp 1666464484
transform 1 0 160608 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1486
timestamp 1666464484
transform 1 0 167776 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1490
timestamp 1666464484
transform 1 0 168224 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_1493
timestamp 1666464484
transform 1 0 168560 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_1557
timestamp 1666464484
transform 1 0 175728 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1561
timestamp 1666464484
transform 1 0 176176 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_129_1564
timestamp 1666464484
transform 1 0 176512 0 -1 105056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1580
timestamp 1666464484
transform 1 0 178304 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_130_2
timestamp 1666464484
transform 1 0 1568 0 1 105056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_34
timestamp 1666464484
transform 1 0 5152 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_37
timestamp 1666464484
transform 1 0 5488 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_101
timestamp 1666464484
transform 1 0 12656 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_105
timestamp 1666464484
transform 1 0 13104 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_108
timestamp 1666464484
transform 1 0 13440 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_172
timestamp 1666464484
transform 1 0 20608 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_176
timestamp 1666464484
transform 1 0 21056 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_179
timestamp 1666464484
transform 1 0 21392 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_243
timestamp 1666464484
transform 1 0 28560 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_247
timestamp 1666464484
transform 1 0 29008 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_250
timestamp 1666464484
transform 1 0 29344 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_314
timestamp 1666464484
transform 1 0 36512 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_318
timestamp 1666464484
transform 1 0 36960 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_321
timestamp 1666464484
transform 1 0 37296 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_385
timestamp 1666464484
transform 1 0 44464 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_389
timestamp 1666464484
transform 1 0 44912 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_392
timestamp 1666464484
transform 1 0 45248 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_456
timestamp 1666464484
transform 1 0 52416 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_460
timestamp 1666464484
transform 1 0 52864 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_463
timestamp 1666464484
transform 1 0 53200 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_527
timestamp 1666464484
transform 1 0 60368 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_531
timestamp 1666464484
transform 1 0 60816 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_534
timestamp 1666464484
transform 1 0 61152 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_598
timestamp 1666464484
transform 1 0 68320 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_602
timestamp 1666464484
transform 1 0 68768 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_605
timestamp 1666464484
transform 1 0 69104 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_669
timestamp 1666464484
transform 1 0 76272 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_673
timestamp 1666464484
transform 1 0 76720 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_676
timestamp 1666464484
transform 1 0 77056 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_740
timestamp 1666464484
transform 1 0 84224 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_744
timestamp 1666464484
transform 1 0 84672 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_747
timestamp 1666464484
transform 1 0 85008 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_811
timestamp 1666464484
transform 1 0 92176 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_815
timestamp 1666464484
transform 1 0 92624 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_818
timestamp 1666464484
transform 1 0 92960 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_882
timestamp 1666464484
transform 1 0 100128 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_886
timestamp 1666464484
transform 1 0 100576 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_889
timestamp 1666464484
transform 1 0 100912 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_953
timestamp 1666464484
transform 1 0 108080 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_957
timestamp 1666464484
transform 1 0 108528 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_960
timestamp 1666464484
transform 1 0 108864 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1024
timestamp 1666464484
transform 1 0 116032 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1028
timestamp 1666464484
transform 1 0 116480 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_1031
timestamp 1666464484
transform 1 0 116816 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1095
timestamp 1666464484
transform 1 0 123984 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1099
timestamp 1666464484
transform 1 0 124432 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_1102
timestamp 1666464484
transform 1 0 124768 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1166
timestamp 1666464484
transform 1 0 131936 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1170
timestamp 1666464484
transform 1 0 132384 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_1173
timestamp 1666464484
transform 1 0 132720 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1237
timestamp 1666464484
transform 1 0 139888 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1241
timestamp 1666464484
transform 1 0 140336 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_1244
timestamp 1666464484
transform 1 0 140672 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1308
timestamp 1666464484
transform 1 0 147840 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1312
timestamp 1666464484
transform 1 0 148288 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_1315
timestamp 1666464484
transform 1 0 148624 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1379
timestamp 1666464484
transform 1 0 155792 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1383
timestamp 1666464484
transform 1 0 156240 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_1386
timestamp 1666464484
transform 1 0 156576 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1450
timestamp 1666464484
transform 1 0 163744 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1454
timestamp 1666464484
transform 1 0 164192 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_1457
timestamp 1666464484
transform 1 0 164528 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1521
timestamp 1666464484
transform 1 0 171696 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1525
timestamp 1666464484
transform 1 0 172144 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_130_1528
timestamp 1666464484
transform 1 0 172480 0 1 105056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_130_1560
timestamp 1666464484
transform 1 0 176064 0 1 105056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1576
timestamp 1666464484
transform 1 0 177856 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1580
timestamp 1666464484
transform 1 0 178304 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_2
timestamp 1666464484
transform 1 0 1568 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_66
timestamp 1666464484
transform 1 0 8736 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_70
timestamp 1666464484
transform 1 0 9184 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_73
timestamp 1666464484
transform 1 0 9520 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_137
timestamp 1666464484
transform 1 0 16688 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_141
timestamp 1666464484
transform 1 0 17136 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_144
timestamp 1666464484
transform 1 0 17472 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_208
timestamp 1666464484
transform 1 0 24640 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_212
timestamp 1666464484
transform 1 0 25088 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_215
timestamp 1666464484
transform 1 0 25424 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_279
timestamp 1666464484
transform 1 0 32592 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_283
timestamp 1666464484
transform 1 0 33040 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_286
timestamp 1666464484
transform 1 0 33376 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_350
timestamp 1666464484
transform 1 0 40544 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_354
timestamp 1666464484
transform 1 0 40992 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_357
timestamp 1666464484
transform 1 0 41328 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_421
timestamp 1666464484
transform 1 0 48496 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_425
timestamp 1666464484
transform 1 0 48944 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_428
timestamp 1666464484
transform 1 0 49280 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_492
timestamp 1666464484
transform 1 0 56448 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_496
timestamp 1666464484
transform 1 0 56896 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_499
timestamp 1666464484
transform 1 0 57232 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_563
timestamp 1666464484
transform 1 0 64400 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_567
timestamp 1666464484
transform 1 0 64848 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_570
timestamp 1666464484
transform 1 0 65184 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_634
timestamp 1666464484
transform 1 0 72352 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_638
timestamp 1666464484
transform 1 0 72800 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_641
timestamp 1666464484
transform 1 0 73136 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_705
timestamp 1666464484
transform 1 0 80304 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_709
timestamp 1666464484
transform 1 0 80752 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_712
timestamp 1666464484
transform 1 0 81088 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_776
timestamp 1666464484
transform 1 0 88256 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_780
timestamp 1666464484
transform 1 0 88704 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_783
timestamp 1666464484
transform 1 0 89040 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_847
timestamp 1666464484
transform 1 0 96208 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_851
timestamp 1666464484
transform 1 0 96656 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_854
timestamp 1666464484
transform 1 0 96992 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_918
timestamp 1666464484
transform 1 0 104160 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_922
timestamp 1666464484
transform 1 0 104608 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_925
timestamp 1666464484
transform 1 0 104944 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_989
timestamp 1666464484
transform 1 0 112112 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_993
timestamp 1666464484
transform 1 0 112560 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_996
timestamp 1666464484
transform 1 0 112896 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1060
timestamp 1666464484
transform 1 0 120064 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1064
timestamp 1666464484
transform 1 0 120512 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_1067
timestamp 1666464484
transform 1 0 120848 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1131
timestamp 1666464484
transform 1 0 128016 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1135
timestamp 1666464484
transform 1 0 128464 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_1138
timestamp 1666464484
transform 1 0 128800 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1202
timestamp 1666464484
transform 1 0 135968 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1206
timestamp 1666464484
transform 1 0 136416 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_1209
timestamp 1666464484
transform 1 0 136752 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1273
timestamp 1666464484
transform 1 0 143920 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1277
timestamp 1666464484
transform 1 0 144368 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_1280
timestamp 1666464484
transform 1 0 144704 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1344
timestamp 1666464484
transform 1 0 151872 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1348
timestamp 1666464484
transform 1 0 152320 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_1351
timestamp 1666464484
transform 1 0 152656 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1415
timestamp 1666464484
transform 1 0 159824 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1419
timestamp 1666464484
transform 1 0 160272 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_1422
timestamp 1666464484
transform 1 0 160608 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1486
timestamp 1666464484
transform 1 0 167776 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1490
timestamp 1666464484
transform 1 0 168224 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_1493
timestamp 1666464484
transform 1 0 168560 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_1557
timestamp 1666464484
transform 1 0 175728 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1561
timestamp 1666464484
transform 1 0 176176 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_131_1564
timestamp 1666464484
transform 1 0 176512 0 -1 106624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1580
timestamp 1666464484
transform 1 0 178304 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_132_2
timestamp 1666464484
transform 1 0 1568 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_34
timestamp 1666464484
transform 1 0 5152 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_37
timestamp 1666464484
transform 1 0 5488 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_101
timestamp 1666464484
transform 1 0 12656 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_105
timestamp 1666464484
transform 1 0 13104 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_108
timestamp 1666464484
transform 1 0 13440 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_172
timestamp 1666464484
transform 1 0 20608 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_176
timestamp 1666464484
transform 1 0 21056 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_179
timestamp 1666464484
transform 1 0 21392 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_243
timestamp 1666464484
transform 1 0 28560 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_247
timestamp 1666464484
transform 1 0 29008 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_250
timestamp 1666464484
transform 1 0 29344 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_314
timestamp 1666464484
transform 1 0 36512 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_318
timestamp 1666464484
transform 1 0 36960 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_321
timestamp 1666464484
transform 1 0 37296 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_385
timestamp 1666464484
transform 1 0 44464 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_389
timestamp 1666464484
transform 1 0 44912 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_392
timestamp 1666464484
transform 1 0 45248 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_456
timestamp 1666464484
transform 1 0 52416 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_460
timestamp 1666464484
transform 1 0 52864 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_463
timestamp 1666464484
transform 1 0 53200 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_527
timestamp 1666464484
transform 1 0 60368 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_531
timestamp 1666464484
transform 1 0 60816 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_534
timestamp 1666464484
transform 1 0 61152 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_598
timestamp 1666464484
transform 1 0 68320 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_602
timestamp 1666464484
transform 1 0 68768 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_605
timestamp 1666464484
transform 1 0 69104 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_669
timestamp 1666464484
transform 1 0 76272 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_673
timestamp 1666464484
transform 1 0 76720 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_676
timestamp 1666464484
transform 1 0 77056 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_740
timestamp 1666464484
transform 1 0 84224 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_744
timestamp 1666464484
transform 1 0 84672 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_747
timestamp 1666464484
transform 1 0 85008 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_811
timestamp 1666464484
transform 1 0 92176 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_815
timestamp 1666464484
transform 1 0 92624 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_818
timestamp 1666464484
transform 1 0 92960 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_882
timestamp 1666464484
transform 1 0 100128 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_886
timestamp 1666464484
transform 1 0 100576 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_889
timestamp 1666464484
transform 1 0 100912 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_953
timestamp 1666464484
transform 1 0 108080 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_957
timestamp 1666464484
transform 1 0 108528 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_960
timestamp 1666464484
transform 1 0 108864 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1024
timestamp 1666464484
transform 1 0 116032 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1028
timestamp 1666464484
transform 1 0 116480 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_1031
timestamp 1666464484
transform 1 0 116816 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1095
timestamp 1666464484
transform 1 0 123984 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1099
timestamp 1666464484
transform 1 0 124432 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_1102
timestamp 1666464484
transform 1 0 124768 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1166
timestamp 1666464484
transform 1 0 131936 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1170
timestamp 1666464484
transform 1 0 132384 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_1173
timestamp 1666464484
transform 1 0 132720 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1237
timestamp 1666464484
transform 1 0 139888 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1241
timestamp 1666464484
transform 1 0 140336 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_1244
timestamp 1666464484
transform 1 0 140672 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1308
timestamp 1666464484
transform 1 0 147840 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1312
timestamp 1666464484
transform 1 0 148288 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_1315
timestamp 1666464484
transform 1 0 148624 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1379
timestamp 1666464484
transform 1 0 155792 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1383
timestamp 1666464484
transform 1 0 156240 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_1386
timestamp 1666464484
transform 1 0 156576 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1450
timestamp 1666464484
transform 1 0 163744 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1454
timestamp 1666464484
transform 1 0 164192 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_1457
timestamp 1666464484
transform 1 0 164528 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1521
timestamp 1666464484
transform 1 0 171696 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1525
timestamp 1666464484
transform 1 0 172144 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_132_1528
timestamp 1666464484
transform 1 0 172480 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_132_1560
timestamp 1666464484
transform 1 0 176064 0 1 106624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1576
timestamp 1666464484
transform 1 0 177856 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1580
timestamp 1666464484
transform 1 0 178304 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_2
timestamp 1666464484
transform 1 0 1568 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_66
timestamp 1666464484
transform 1 0 8736 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_70
timestamp 1666464484
transform 1 0 9184 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_73
timestamp 1666464484
transform 1 0 9520 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_137
timestamp 1666464484
transform 1 0 16688 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_141
timestamp 1666464484
transform 1 0 17136 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_144
timestamp 1666464484
transform 1 0 17472 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_208
timestamp 1666464484
transform 1 0 24640 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_212
timestamp 1666464484
transform 1 0 25088 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_215
timestamp 1666464484
transform 1 0 25424 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_279
timestamp 1666464484
transform 1 0 32592 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_283
timestamp 1666464484
transform 1 0 33040 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_286
timestamp 1666464484
transform 1 0 33376 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_350
timestamp 1666464484
transform 1 0 40544 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_354
timestamp 1666464484
transform 1 0 40992 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_357
timestamp 1666464484
transform 1 0 41328 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_421
timestamp 1666464484
transform 1 0 48496 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_425
timestamp 1666464484
transform 1 0 48944 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_428
timestamp 1666464484
transform 1 0 49280 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_492
timestamp 1666464484
transform 1 0 56448 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_496
timestamp 1666464484
transform 1 0 56896 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_499
timestamp 1666464484
transform 1 0 57232 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_563
timestamp 1666464484
transform 1 0 64400 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_567
timestamp 1666464484
transform 1 0 64848 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_570
timestamp 1666464484
transform 1 0 65184 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_634
timestamp 1666464484
transform 1 0 72352 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_638
timestamp 1666464484
transform 1 0 72800 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_641
timestamp 1666464484
transform 1 0 73136 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_705
timestamp 1666464484
transform 1 0 80304 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_709
timestamp 1666464484
transform 1 0 80752 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_712
timestamp 1666464484
transform 1 0 81088 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_776
timestamp 1666464484
transform 1 0 88256 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_780
timestamp 1666464484
transform 1 0 88704 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_783
timestamp 1666464484
transform 1 0 89040 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_847
timestamp 1666464484
transform 1 0 96208 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_851
timestamp 1666464484
transform 1 0 96656 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_854
timestamp 1666464484
transform 1 0 96992 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_918
timestamp 1666464484
transform 1 0 104160 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_922
timestamp 1666464484
transform 1 0 104608 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_925
timestamp 1666464484
transform 1 0 104944 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_989
timestamp 1666464484
transform 1 0 112112 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_993
timestamp 1666464484
transform 1 0 112560 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_996
timestamp 1666464484
transform 1 0 112896 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1060
timestamp 1666464484
transform 1 0 120064 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1064
timestamp 1666464484
transform 1 0 120512 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_1067
timestamp 1666464484
transform 1 0 120848 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1131
timestamp 1666464484
transform 1 0 128016 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1135
timestamp 1666464484
transform 1 0 128464 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_1138
timestamp 1666464484
transform 1 0 128800 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1202
timestamp 1666464484
transform 1 0 135968 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1206
timestamp 1666464484
transform 1 0 136416 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_1209
timestamp 1666464484
transform 1 0 136752 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1273
timestamp 1666464484
transform 1 0 143920 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1277
timestamp 1666464484
transform 1 0 144368 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_1280
timestamp 1666464484
transform 1 0 144704 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1344
timestamp 1666464484
transform 1 0 151872 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1348
timestamp 1666464484
transform 1 0 152320 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_1351
timestamp 1666464484
transform 1 0 152656 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1415
timestamp 1666464484
transform 1 0 159824 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1419
timestamp 1666464484
transform 1 0 160272 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_1422
timestamp 1666464484
transform 1 0 160608 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1486
timestamp 1666464484
transform 1 0 167776 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1490
timestamp 1666464484
transform 1 0 168224 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_1493
timestamp 1666464484
transform 1 0 168560 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1557
timestamp 1666464484
transform 1 0 175728 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1561
timestamp 1666464484
transform 1 0 176176 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_133_1564
timestamp 1666464484
transform 1 0 176512 0 -1 108192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1580
timestamp 1666464484
transform 1 0 178304 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_134_2
timestamp 1666464484
transform 1 0 1568 0 1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_34
timestamp 1666464484
transform 1 0 5152 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_37
timestamp 1666464484
transform 1 0 5488 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_101
timestamp 1666464484
transform 1 0 12656 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_105
timestamp 1666464484
transform 1 0 13104 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_108
timestamp 1666464484
transform 1 0 13440 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_172
timestamp 1666464484
transform 1 0 20608 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_176
timestamp 1666464484
transform 1 0 21056 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_179
timestamp 1666464484
transform 1 0 21392 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_243
timestamp 1666464484
transform 1 0 28560 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_247
timestamp 1666464484
transform 1 0 29008 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_250
timestamp 1666464484
transform 1 0 29344 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_314
timestamp 1666464484
transform 1 0 36512 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_318
timestamp 1666464484
transform 1 0 36960 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_321
timestamp 1666464484
transform 1 0 37296 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_385
timestamp 1666464484
transform 1 0 44464 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_389
timestamp 1666464484
transform 1 0 44912 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_392
timestamp 1666464484
transform 1 0 45248 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_456
timestamp 1666464484
transform 1 0 52416 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_460
timestamp 1666464484
transform 1 0 52864 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_463
timestamp 1666464484
transform 1 0 53200 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_527
timestamp 1666464484
transform 1 0 60368 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_531
timestamp 1666464484
transform 1 0 60816 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_534
timestamp 1666464484
transform 1 0 61152 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_598
timestamp 1666464484
transform 1 0 68320 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_602
timestamp 1666464484
transform 1 0 68768 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_605
timestamp 1666464484
transform 1 0 69104 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_669
timestamp 1666464484
transform 1 0 76272 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_673
timestamp 1666464484
transform 1 0 76720 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_676
timestamp 1666464484
transform 1 0 77056 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_740
timestamp 1666464484
transform 1 0 84224 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_744
timestamp 1666464484
transform 1 0 84672 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_747
timestamp 1666464484
transform 1 0 85008 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_811
timestamp 1666464484
transform 1 0 92176 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_815
timestamp 1666464484
transform 1 0 92624 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_818
timestamp 1666464484
transform 1 0 92960 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_882
timestamp 1666464484
transform 1 0 100128 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_886
timestamp 1666464484
transform 1 0 100576 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_889
timestamp 1666464484
transform 1 0 100912 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_953
timestamp 1666464484
transform 1 0 108080 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_957
timestamp 1666464484
transform 1 0 108528 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_960
timestamp 1666464484
transform 1 0 108864 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1024
timestamp 1666464484
transform 1 0 116032 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1028
timestamp 1666464484
transform 1 0 116480 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_1031
timestamp 1666464484
transform 1 0 116816 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1095
timestamp 1666464484
transform 1 0 123984 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1099
timestamp 1666464484
transform 1 0 124432 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_1102
timestamp 1666464484
transform 1 0 124768 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1166
timestamp 1666464484
transform 1 0 131936 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1170
timestamp 1666464484
transform 1 0 132384 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_1173
timestamp 1666464484
transform 1 0 132720 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1237
timestamp 1666464484
transform 1 0 139888 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1241
timestamp 1666464484
transform 1 0 140336 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_1244
timestamp 1666464484
transform 1 0 140672 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1308
timestamp 1666464484
transform 1 0 147840 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1312
timestamp 1666464484
transform 1 0 148288 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_1315
timestamp 1666464484
transform 1 0 148624 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1379
timestamp 1666464484
transform 1 0 155792 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1383
timestamp 1666464484
transform 1 0 156240 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_1386
timestamp 1666464484
transform 1 0 156576 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1450
timestamp 1666464484
transform 1 0 163744 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1454
timestamp 1666464484
transform 1 0 164192 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_1457
timestamp 1666464484
transform 1 0 164528 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1521
timestamp 1666464484
transform 1 0 171696 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1525
timestamp 1666464484
transform 1 0 172144 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_134_1528
timestamp 1666464484
transform 1 0 172480 0 1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_134_1560
timestamp 1666464484
transform 1 0 176064 0 1 108192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1576
timestamp 1666464484
transform 1 0 177856 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1580
timestamp 1666464484
transform 1 0 178304 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_2
timestamp 1666464484
transform 1 0 1568 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_66
timestamp 1666464484
transform 1 0 8736 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_70
timestamp 1666464484
transform 1 0 9184 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_73
timestamp 1666464484
transform 1 0 9520 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_137
timestamp 1666464484
transform 1 0 16688 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_141
timestamp 1666464484
transform 1 0 17136 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_144
timestamp 1666464484
transform 1 0 17472 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_208
timestamp 1666464484
transform 1 0 24640 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_212
timestamp 1666464484
transform 1 0 25088 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_215
timestamp 1666464484
transform 1 0 25424 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_279
timestamp 1666464484
transform 1 0 32592 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_283
timestamp 1666464484
transform 1 0 33040 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_286
timestamp 1666464484
transform 1 0 33376 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_350
timestamp 1666464484
transform 1 0 40544 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_354
timestamp 1666464484
transform 1 0 40992 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_357
timestamp 1666464484
transform 1 0 41328 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_421
timestamp 1666464484
transform 1 0 48496 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_425
timestamp 1666464484
transform 1 0 48944 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_428
timestamp 1666464484
transform 1 0 49280 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_492
timestamp 1666464484
transform 1 0 56448 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_496
timestamp 1666464484
transform 1 0 56896 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_499
timestamp 1666464484
transform 1 0 57232 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_563
timestamp 1666464484
transform 1 0 64400 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_567
timestamp 1666464484
transform 1 0 64848 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_570
timestamp 1666464484
transform 1 0 65184 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_634
timestamp 1666464484
transform 1 0 72352 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_638
timestamp 1666464484
transform 1 0 72800 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_641
timestamp 1666464484
transform 1 0 73136 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_705
timestamp 1666464484
transform 1 0 80304 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_709
timestamp 1666464484
transform 1 0 80752 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_712
timestamp 1666464484
transform 1 0 81088 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_776
timestamp 1666464484
transform 1 0 88256 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_780
timestamp 1666464484
transform 1 0 88704 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_783
timestamp 1666464484
transform 1 0 89040 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_847
timestamp 1666464484
transform 1 0 96208 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_851
timestamp 1666464484
transform 1 0 96656 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_854
timestamp 1666464484
transform 1 0 96992 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_918
timestamp 1666464484
transform 1 0 104160 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_922
timestamp 1666464484
transform 1 0 104608 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_925
timestamp 1666464484
transform 1 0 104944 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_989
timestamp 1666464484
transform 1 0 112112 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_993
timestamp 1666464484
transform 1 0 112560 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_996
timestamp 1666464484
transform 1 0 112896 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1060
timestamp 1666464484
transform 1 0 120064 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1064
timestamp 1666464484
transform 1 0 120512 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_1067
timestamp 1666464484
transform 1 0 120848 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1131
timestamp 1666464484
transform 1 0 128016 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1135
timestamp 1666464484
transform 1 0 128464 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_1138
timestamp 1666464484
transform 1 0 128800 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1202
timestamp 1666464484
transform 1 0 135968 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1206
timestamp 1666464484
transform 1 0 136416 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_1209
timestamp 1666464484
transform 1 0 136752 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1273
timestamp 1666464484
transform 1 0 143920 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1277
timestamp 1666464484
transform 1 0 144368 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_1280
timestamp 1666464484
transform 1 0 144704 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1344
timestamp 1666464484
transform 1 0 151872 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1348
timestamp 1666464484
transform 1 0 152320 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_1351
timestamp 1666464484
transform 1 0 152656 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1415
timestamp 1666464484
transform 1 0 159824 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1419
timestamp 1666464484
transform 1 0 160272 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_1422
timestamp 1666464484
transform 1 0 160608 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1486
timestamp 1666464484
transform 1 0 167776 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1490
timestamp 1666464484
transform 1 0 168224 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_1493
timestamp 1666464484
transform 1 0 168560 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_1557
timestamp 1666464484
transform 1 0 175728 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1561
timestamp 1666464484
transform 1 0 176176 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_135_1564
timestamp 1666464484
transform 1 0 176512 0 -1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1580
timestamp 1666464484
transform 1 0 178304 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_136_2
timestamp 1666464484
transform 1 0 1568 0 1 109760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_34
timestamp 1666464484
transform 1 0 5152 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_37
timestamp 1666464484
transform 1 0 5488 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_101
timestamp 1666464484
transform 1 0 12656 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_105
timestamp 1666464484
transform 1 0 13104 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_108
timestamp 1666464484
transform 1 0 13440 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_172
timestamp 1666464484
transform 1 0 20608 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_176
timestamp 1666464484
transform 1 0 21056 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_179
timestamp 1666464484
transform 1 0 21392 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_243
timestamp 1666464484
transform 1 0 28560 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_247
timestamp 1666464484
transform 1 0 29008 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_250
timestamp 1666464484
transform 1 0 29344 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_314
timestamp 1666464484
transform 1 0 36512 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_318
timestamp 1666464484
transform 1 0 36960 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_321
timestamp 1666464484
transform 1 0 37296 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_385
timestamp 1666464484
transform 1 0 44464 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_389
timestamp 1666464484
transform 1 0 44912 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_392
timestamp 1666464484
transform 1 0 45248 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_456
timestamp 1666464484
transform 1 0 52416 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_460
timestamp 1666464484
transform 1 0 52864 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_463
timestamp 1666464484
transform 1 0 53200 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_527
timestamp 1666464484
transform 1 0 60368 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_531
timestamp 1666464484
transform 1 0 60816 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_534
timestamp 1666464484
transform 1 0 61152 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_598
timestamp 1666464484
transform 1 0 68320 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_602
timestamp 1666464484
transform 1 0 68768 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_605
timestamp 1666464484
transform 1 0 69104 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_669
timestamp 1666464484
transform 1 0 76272 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_673
timestamp 1666464484
transform 1 0 76720 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_676
timestamp 1666464484
transform 1 0 77056 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_740
timestamp 1666464484
transform 1 0 84224 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_744
timestamp 1666464484
transform 1 0 84672 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_747
timestamp 1666464484
transform 1 0 85008 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_811
timestamp 1666464484
transform 1 0 92176 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_815
timestamp 1666464484
transform 1 0 92624 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_818
timestamp 1666464484
transform 1 0 92960 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_882
timestamp 1666464484
transform 1 0 100128 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_886
timestamp 1666464484
transform 1 0 100576 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_889
timestamp 1666464484
transform 1 0 100912 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_953
timestamp 1666464484
transform 1 0 108080 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_957
timestamp 1666464484
transform 1 0 108528 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_960
timestamp 1666464484
transform 1 0 108864 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1024
timestamp 1666464484
transform 1 0 116032 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1028
timestamp 1666464484
transform 1 0 116480 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_1031
timestamp 1666464484
transform 1 0 116816 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1095
timestamp 1666464484
transform 1 0 123984 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1099
timestamp 1666464484
transform 1 0 124432 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_1102
timestamp 1666464484
transform 1 0 124768 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1166
timestamp 1666464484
transform 1 0 131936 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1170
timestamp 1666464484
transform 1 0 132384 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_1173
timestamp 1666464484
transform 1 0 132720 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1237
timestamp 1666464484
transform 1 0 139888 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1241
timestamp 1666464484
transform 1 0 140336 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_1244
timestamp 1666464484
transform 1 0 140672 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1308
timestamp 1666464484
transform 1 0 147840 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1312
timestamp 1666464484
transform 1 0 148288 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_1315
timestamp 1666464484
transform 1 0 148624 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1379
timestamp 1666464484
transform 1 0 155792 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1383
timestamp 1666464484
transform 1 0 156240 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_1386
timestamp 1666464484
transform 1 0 156576 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1450
timestamp 1666464484
transform 1 0 163744 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1454
timestamp 1666464484
transform 1 0 164192 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_1457
timestamp 1666464484
transform 1 0 164528 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1521
timestamp 1666464484
transform 1 0 171696 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1525
timestamp 1666464484
transform 1 0 172144 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_136_1528
timestamp 1666464484
transform 1 0 172480 0 1 109760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_136_1560
timestamp 1666464484
transform 1 0 176064 0 1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1576
timestamp 1666464484
transform 1 0 177856 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1580
timestamp 1666464484
transform 1 0 178304 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_2
timestamp 1666464484
transform 1 0 1568 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_66
timestamp 1666464484
transform 1 0 8736 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_70
timestamp 1666464484
transform 1 0 9184 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_73
timestamp 1666464484
transform 1 0 9520 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_137
timestamp 1666464484
transform 1 0 16688 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_141
timestamp 1666464484
transform 1 0 17136 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_144
timestamp 1666464484
transform 1 0 17472 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_208
timestamp 1666464484
transform 1 0 24640 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_212
timestamp 1666464484
transform 1 0 25088 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_215
timestamp 1666464484
transform 1 0 25424 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_279
timestamp 1666464484
transform 1 0 32592 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_283
timestamp 1666464484
transform 1 0 33040 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_286
timestamp 1666464484
transform 1 0 33376 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_350
timestamp 1666464484
transform 1 0 40544 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_354
timestamp 1666464484
transform 1 0 40992 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_357
timestamp 1666464484
transform 1 0 41328 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_421
timestamp 1666464484
transform 1 0 48496 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_425
timestamp 1666464484
transform 1 0 48944 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_428
timestamp 1666464484
transform 1 0 49280 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_492
timestamp 1666464484
transform 1 0 56448 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_496
timestamp 1666464484
transform 1 0 56896 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_499
timestamp 1666464484
transform 1 0 57232 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_563
timestamp 1666464484
transform 1 0 64400 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_567
timestamp 1666464484
transform 1 0 64848 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_570
timestamp 1666464484
transform 1 0 65184 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_634
timestamp 1666464484
transform 1 0 72352 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_638
timestamp 1666464484
transform 1 0 72800 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_641
timestamp 1666464484
transform 1 0 73136 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_705
timestamp 1666464484
transform 1 0 80304 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_709
timestamp 1666464484
transform 1 0 80752 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_712
timestamp 1666464484
transform 1 0 81088 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_776
timestamp 1666464484
transform 1 0 88256 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_780
timestamp 1666464484
transform 1 0 88704 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_783
timestamp 1666464484
transform 1 0 89040 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_847
timestamp 1666464484
transform 1 0 96208 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_851
timestamp 1666464484
transform 1 0 96656 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_854
timestamp 1666464484
transform 1 0 96992 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_918
timestamp 1666464484
transform 1 0 104160 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_922
timestamp 1666464484
transform 1 0 104608 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_925
timestamp 1666464484
transform 1 0 104944 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_989
timestamp 1666464484
transform 1 0 112112 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_993
timestamp 1666464484
transform 1 0 112560 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_996
timestamp 1666464484
transform 1 0 112896 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1060
timestamp 1666464484
transform 1 0 120064 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1064
timestamp 1666464484
transform 1 0 120512 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_1067
timestamp 1666464484
transform 1 0 120848 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1131
timestamp 1666464484
transform 1 0 128016 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1135
timestamp 1666464484
transform 1 0 128464 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_1138
timestamp 1666464484
transform 1 0 128800 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1202
timestamp 1666464484
transform 1 0 135968 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1206
timestamp 1666464484
transform 1 0 136416 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_1209
timestamp 1666464484
transform 1 0 136752 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1273
timestamp 1666464484
transform 1 0 143920 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1277
timestamp 1666464484
transform 1 0 144368 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_1280
timestamp 1666464484
transform 1 0 144704 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1344
timestamp 1666464484
transform 1 0 151872 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1348
timestamp 1666464484
transform 1 0 152320 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_1351
timestamp 1666464484
transform 1 0 152656 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1415
timestamp 1666464484
transform 1 0 159824 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1419
timestamp 1666464484
transform 1 0 160272 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_1422
timestamp 1666464484
transform 1 0 160608 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1486
timestamp 1666464484
transform 1 0 167776 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1490
timestamp 1666464484
transform 1 0 168224 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_1493
timestamp 1666464484
transform 1 0 168560 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1557
timestamp 1666464484
transform 1 0 175728 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1561
timestamp 1666464484
transform 1 0 176176 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_137_1564
timestamp 1666464484
transform 1 0 176512 0 -1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1580
timestamp 1666464484
transform 1 0 178304 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_138_2
timestamp 1666464484
transform 1 0 1568 0 1 111328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_34
timestamp 1666464484
transform 1 0 5152 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_37
timestamp 1666464484
transform 1 0 5488 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_101
timestamp 1666464484
transform 1 0 12656 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_105
timestamp 1666464484
transform 1 0 13104 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_108
timestamp 1666464484
transform 1 0 13440 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_172
timestamp 1666464484
transform 1 0 20608 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_176
timestamp 1666464484
transform 1 0 21056 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_179
timestamp 1666464484
transform 1 0 21392 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_243
timestamp 1666464484
transform 1 0 28560 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_247
timestamp 1666464484
transform 1 0 29008 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_250
timestamp 1666464484
transform 1 0 29344 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_314
timestamp 1666464484
transform 1 0 36512 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_318
timestamp 1666464484
transform 1 0 36960 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_321
timestamp 1666464484
transform 1 0 37296 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_385
timestamp 1666464484
transform 1 0 44464 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_389
timestamp 1666464484
transform 1 0 44912 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_392
timestamp 1666464484
transform 1 0 45248 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_456
timestamp 1666464484
transform 1 0 52416 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_460
timestamp 1666464484
transform 1 0 52864 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_463
timestamp 1666464484
transform 1 0 53200 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_527
timestamp 1666464484
transform 1 0 60368 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_531
timestamp 1666464484
transform 1 0 60816 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_534
timestamp 1666464484
transform 1 0 61152 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_598
timestamp 1666464484
transform 1 0 68320 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_602
timestamp 1666464484
transform 1 0 68768 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_605
timestamp 1666464484
transform 1 0 69104 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_669
timestamp 1666464484
transform 1 0 76272 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_673
timestamp 1666464484
transform 1 0 76720 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_676
timestamp 1666464484
transform 1 0 77056 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_740
timestamp 1666464484
transform 1 0 84224 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_744
timestamp 1666464484
transform 1 0 84672 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_747
timestamp 1666464484
transform 1 0 85008 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_811
timestamp 1666464484
transform 1 0 92176 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_815
timestamp 1666464484
transform 1 0 92624 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_818
timestamp 1666464484
transform 1 0 92960 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_882
timestamp 1666464484
transform 1 0 100128 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_886
timestamp 1666464484
transform 1 0 100576 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_889
timestamp 1666464484
transform 1 0 100912 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_953
timestamp 1666464484
transform 1 0 108080 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_957
timestamp 1666464484
transform 1 0 108528 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_960
timestamp 1666464484
transform 1 0 108864 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1024
timestamp 1666464484
transform 1 0 116032 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1028
timestamp 1666464484
transform 1 0 116480 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_1031
timestamp 1666464484
transform 1 0 116816 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1095
timestamp 1666464484
transform 1 0 123984 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1099
timestamp 1666464484
transform 1 0 124432 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_1102
timestamp 1666464484
transform 1 0 124768 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1166
timestamp 1666464484
transform 1 0 131936 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1170
timestamp 1666464484
transform 1 0 132384 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_1173
timestamp 1666464484
transform 1 0 132720 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1237
timestamp 1666464484
transform 1 0 139888 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1241
timestamp 1666464484
transform 1 0 140336 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_1244
timestamp 1666464484
transform 1 0 140672 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1308
timestamp 1666464484
transform 1 0 147840 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1312
timestamp 1666464484
transform 1 0 148288 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_1315
timestamp 1666464484
transform 1 0 148624 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1379
timestamp 1666464484
transform 1 0 155792 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1383
timestamp 1666464484
transform 1 0 156240 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_1386
timestamp 1666464484
transform 1 0 156576 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1450
timestamp 1666464484
transform 1 0 163744 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1454
timestamp 1666464484
transform 1 0 164192 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_1457
timestamp 1666464484
transform 1 0 164528 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1521
timestamp 1666464484
transform 1 0 171696 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1525
timestamp 1666464484
transform 1 0 172144 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_138_1528
timestamp 1666464484
transform 1 0 172480 0 1 111328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_138_1560
timestamp 1666464484
transform 1 0 176064 0 1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1576
timestamp 1666464484
transform 1 0 177856 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1580
timestamp 1666464484
transform 1 0 178304 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_2
timestamp 1666464484
transform 1 0 1568 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_66
timestamp 1666464484
transform 1 0 8736 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_70
timestamp 1666464484
transform 1 0 9184 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_73
timestamp 1666464484
transform 1 0 9520 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_137
timestamp 1666464484
transform 1 0 16688 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_141
timestamp 1666464484
transform 1 0 17136 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_144
timestamp 1666464484
transform 1 0 17472 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_208
timestamp 1666464484
transform 1 0 24640 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_212
timestamp 1666464484
transform 1 0 25088 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_215
timestamp 1666464484
transform 1 0 25424 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_279
timestamp 1666464484
transform 1 0 32592 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_283
timestamp 1666464484
transform 1 0 33040 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_286
timestamp 1666464484
transform 1 0 33376 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_350
timestamp 1666464484
transform 1 0 40544 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_354
timestamp 1666464484
transform 1 0 40992 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_357
timestamp 1666464484
transform 1 0 41328 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_421
timestamp 1666464484
transform 1 0 48496 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_425
timestamp 1666464484
transform 1 0 48944 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_428
timestamp 1666464484
transform 1 0 49280 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_492
timestamp 1666464484
transform 1 0 56448 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_496
timestamp 1666464484
transform 1 0 56896 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_499
timestamp 1666464484
transform 1 0 57232 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_563
timestamp 1666464484
transform 1 0 64400 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_567
timestamp 1666464484
transform 1 0 64848 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_570
timestamp 1666464484
transform 1 0 65184 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_634
timestamp 1666464484
transform 1 0 72352 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_638
timestamp 1666464484
transform 1 0 72800 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_641
timestamp 1666464484
transform 1 0 73136 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_705
timestamp 1666464484
transform 1 0 80304 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_709
timestamp 1666464484
transform 1 0 80752 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_712
timestamp 1666464484
transform 1 0 81088 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_776
timestamp 1666464484
transform 1 0 88256 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_780
timestamp 1666464484
transform 1 0 88704 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_783
timestamp 1666464484
transform 1 0 89040 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_847
timestamp 1666464484
transform 1 0 96208 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_851
timestamp 1666464484
transform 1 0 96656 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_854
timestamp 1666464484
transform 1 0 96992 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_918
timestamp 1666464484
transform 1 0 104160 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_922
timestamp 1666464484
transform 1 0 104608 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_925
timestamp 1666464484
transform 1 0 104944 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_989
timestamp 1666464484
transform 1 0 112112 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_993
timestamp 1666464484
transform 1 0 112560 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_996
timestamp 1666464484
transform 1 0 112896 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1060
timestamp 1666464484
transform 1 0 120064 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1064
timestamp 1666464484
transform 1 0 120512 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_1067
timestamp 1666464484
transform 1 0 120848 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1131
timestamp 1666464484
transform 1 0 128016 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1135
timestamp 1666464484
transform 1 0 128464 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_1138
timestamp 1666464484
transform 1 0 128800 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1202
timestamp 1666464484
transform 1 0 135968 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1206
timestamp 1666464484
transform 1 0 136416 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_1209
timestamp 1666464484
transform 1 0 136752 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1273
timestamp 1666464484
transform 1 0 143920 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1277
timestamp 1666464484
transform 1 0 144368 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_1280
timestamp 1666464484
transform 1 0 144704 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1344
timestamp 1666464484
transform 1 0 151872 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1348
timestamp 1666464484
transform 1 0 152320 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_1351
timestamp 1666464484
transform 1 0 152656 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1415
timestamp 1666464484
transform 1 0 159824 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1419
timestamp 1666464484
transform 1 0 160272 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_1422
timestamp 1666464484
transform 1 0 160608 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1486
timestamp 1666464484
transform 1 0 167776 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1490
timestamp 1666464484
transform 1 0 168224 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_1493
timestamp 1666464484
transform 1 0 168560 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_1557
timestamp 1666464484
transform 1 0 175728 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1561
timestamp 1666464484
transform 1 0 176176 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_139_1564
timestamp 1666464484
transform 1 0 176512 0 -1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1580
timestamp 1666464484
transform 1 0 178304 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_140_2
timestamp 1666464484
transform 1 0 1568 0 1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_34
timestamp 1666464484
transform 1 0 5152 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_37
timestamp 1666464484
transform 1 0 5488 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_101
timestamp 1666464484
transform 1 0 12656 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_105
timestamp 1666464484
transform 1 0 13104 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_108
timestamp 1666464484
transform 1 0 13440 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_172
timestamp 1666464484
transform 1 0 20608 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_176
timestamp 1666464484
transform 1 0 21056 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_179
timestamp 1666464484
transform 1 0 21392 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_243
timestamp 1666464484
transform 1 0 28560 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_247
timestamp 1666464484
transform 1 0 29008 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_250
timestamp 1666464484
transform 1 0 29344 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_314
timestamp 1666464484
transform 1 0 36512 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_318
timestamp 1666464484
transform 1 0 36960 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_321
timestamp 1666464484
transform 1 0 37296 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_385
timestamp 1666464484
transform 1 0 44464 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_389
timestamp 1666464484
transform 1 0 44912 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_392
timestamp 1666464484
transform 1 0 45248 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_456
timestamp 1666464484
transform 1 0 52416 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_460
timestamp 1666464484
transform 1 0 52864 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_463
timestamp 1666464484
transform 1 0 53200 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_527
timestamp 1666464484
transform 1 0 60368 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_531
timestamp 1666464484
transform 1 0 60816 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_534
timestamp 1666464484
transform 1 0 61152 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_598
timestamp 1666464484
transform 1 0 68320 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_602
timestamp 1666464484
transform 1 0 68768 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_605
timestamp 1666464484
transform 1 0 69104 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_669
timestamp 1666464484
transform 1 0 76272 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_673
timestamp 1666464484
transform 1 0 76720 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_676
timestamp 1666464484
transform 1 0 77056 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_740
timestamp 1666464484
transform 1 0 84224 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_744
timestamp 1666464484
transform 1 0 84672 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_747
timestamp 1666464484
transform 1 0 85008 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_811
timestamp 1666464484
transform 1 0 92176 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_815
timestamp 1666464484
transform 1 0 92624 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_818
timestamp 1666464484
transform 1 0 92960 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_882
timestamp 1666464484
transform 1 0 100128 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_886
timestamp 1666464484
transform 1 0 100576 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_889
timestamp 1666464484
transform 1 0 100912 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_953
timestamp 1666464484
transform 1 0 108080 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_957
timestamp 1666464484
transform 1 0 108528 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_960
timestamp 1666464484
transform 1 0 108864 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1024
timestamp 1666464484
transform 1 0 116032 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1028
timestamp 1666464484
transform 1 0 116480 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_1031
timestamp 1666464484
transform 1 0 116816 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1095
timestamp 1666464484
transform 1 0 123984 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1099
timestamp 1666464484
transform 1 0 124432 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_1102
timestamp 1666464484
transform 1 0 124768 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1166
timestamp 1666464484
transform 1 0 131936 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1170
timestamp 1666464484
transform 1 0 132384 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_1173
timestamp 1666464484
transform 1 0 132720 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1237
timestamp 1666464484
transform 1 0 139888 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1241
timestamp 1666464484
transform 1 0 140336 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_1244
timestamp 1666464484
transform 1 0 140672 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1308
timestamp 1666464484
transform 1 0 147840 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1312
timestamp 1666464484
transform 1 0 148288 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_1315
timestamp 1666464484
transform 1 0 148624 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1379
timestamp 1666464484
transform 1 0 155792 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1383
timestamp 1666464484
transform 1 0 156240 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_1386
timestamp 1666464484
transform 1 0 156576 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1450
timestamp 1666464484
transform 1 0 163744 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1454
timestamp 1666464484
transform 1 0 164192 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_1457
timestamp 1666464484
transform 1 0 164528 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1521
timestamp 1666464484
transform 1 0 171696 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1525
timestamp 1666464484
transform 1 0 172144 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_140_1528
timestamp 1666464484
transform 1 0 172480 0 1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_140_1560
timestamp 1666464484
transform 1 0 176064 0 1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1576
timestamp 1666464484
transform 1 0 177856 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1580
timestamp 1666464484
transform 1 0 178304 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_2
timestamp 1666464484
transform 1 0 1568 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_66
timestamp 1666464484
transform 1 0 8736 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_70
timestamp 1666464484
transform 1 0 9184 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_73
timestamp 1666464484
transform 1 0 9520 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_137
timestamp 1666464484
transform 1 0 16688 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_141
timestamp 1666464484
transform 1 0 17136 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_144
timestamp 1666464484
transform 1 0 17472 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_208
timestamp 1666464484
transform 1 0 24640 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_212
timestamp 1666464484
transform 1 0 25088 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_215
timestamp 1666464484
transform 1 0 25424 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_279
timestamp 1666464484
transform 1 0 32592 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_283
timestamp 1666464484
transform 1 0 33040 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_286
timestamp 1666464484
transform 1 0 33376 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_350
timestamp 1666464484
transform 1 0 40544 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_354
timestamp 1666464484
transform 1 0 40992 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_357
timestamp 1666464484
transform 1 0 41328 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_421
timestamp 1666464484
transform 1 0 48496 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_425
timestamp 1666464484
transform 1 0 48944 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_428
timestamp 1666464484
transform 1 0 49280 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_492
timestamp 1666464484
transform 1 0 56448 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_496
timestamp 1666464484
transform 1 0 56896 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_499
timestamp 1666464484
transform 1 0 57232 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_563
timestamp 1666464484
transform 1 0 64400 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_567
timestamp 1666464484
transform 1 0 64848 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_570
timestamp 1666464484
transform 1 0 65184 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_634
timestamp 1666464484
transform 1 0 72352 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_638
timestamp 1666464484
transform 1 0 72800 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_641
timestamp 1666464484
transform 1 0 73136 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_705
timestamp 1666464484
transform 1 0 80304 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_709
timestamp 1666464484
transform 1 0 80752 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_712
timestamp 1666464484
transform 1 0 81088 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_776
timestamp 1666464484
transform 1 0 88256 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_780
timestamp 1666464484
transform 1 0 88704 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_783
timestamp 1666464484
transform 1 0 89040 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_847
timestamp 1666464484
transform 1 0 96208 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_851
timestamp 1666464484
transform 1 0 96656 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_854
timestamp 1666464484
transform 1 0 96992 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_918
timestamp 1666464484
transform 1 0 104160 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_922
timestamp 1666464484
transform 1 0 104608 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_925
timestamp 1666464484
transform 1 0 104944 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_989
timestamp 1666464484
transform 1 0 112112 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_993
timestamp 1666464484
transform 1 0 112560 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_996
timestamp 1666464484
transform 1 0 112896 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1060
timestamp 1666464484
transform 1 0 120064 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1064
timestamp 1666464484
transform 1 0 120512 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_1067
timestamp 1666464484
transform 1 0 120848 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1131
timestamp 1666464484
transform 1 0 128016 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1135
timestamp 1666464484
transform 1 0 128464 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_1138
timestamp 1666464484
transform 1 0 128800 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1202
timestamp 1666464484
transform 1 0 135968 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1206
timestamp 1666464484
transform 1 0 136416 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_1209
timestamp 1666464484
transform 1 0 136752 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1273
timestamp 1666464484
transform 1 0 143920 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1277
timestamp 1666464484
transform 1 0 144368 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_1280
timestamp 1666464484
transform 1 0 144704 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1344
timestamp 1666464484
transform 1 0 151872 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1348
timestamp 1666464484
transform 1 0 152320 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_1351
timestamp 1666464484
transform 1 0 152656 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1415
timestamp 1666464484
transform 1 0 159824 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1419
timestamp 1666464484
transform 1 0 160272 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_1422
timestamp 1666464484
transform 1 0 160608 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1486
timestamp 1666464484
transform 1 0 167776 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1490
timestamp 1666464484
transform 1 0 168224 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_1493
timestamp 1666464484
transform 1 0 168560 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1557
timestamp 1666464484
transform 1 0 175728 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1561
timestamp 1666464484
transform 1 0 176176 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_141_1564
timestamp 1666464484
transform 1 0 176512 0 -1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1580
timestamp 1666464484
transform 1 0 178304 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_2
timestamp 1666464484
transform 1 0 1568 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_34
timestamp 1666464484
transform 1 0 5152 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_37
timestamp 1666464484
transform 1 0 5488 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_101
timestamp 1666464484
transform 1 0 12656 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_105
timestamp 1666464484
transform 1 0 13104 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_108
timestamp 1666464484
transform 1 0 13440 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_172
timestamp 1666464484
transform 1 0 20608 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_176
timestamp 1666464484
transform 1 0 21056 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_179
timestamp 1666464484
transform 1 0 21392 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_243
timestamp 1666464484
transform 1 0 28560 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_247
timestamp 1666464484
transform 1 0 29008 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_250
timestamp 1666464484
transform 1 0 29344 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_314
timestamp 1666464484
transform 1 0 36512 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_318
timestamp 1666464484
transform 1 0 36960 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_321
timestamp 1666464484
transform 1 0 37296 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_385
timestamp 1666464484
transform 1 0 44464 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_389
timestamp 1666464484
transform 1 0 44912 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_392
timestamp 1666464484
transform 1 0 45248 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_456
timestamp 1666464484
transform 1 0 52416 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_460
timestamp 1666464484
transform 1 0 52864 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_463
timestamp 1666464484
transform 1 0 53200 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_527
timestamp 1666464484
transform 1 0 60368 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_531
timestamp 1666464484
transform 1 0 60816 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_534
timestamp 1666464484
transform 1 0 61152 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_550
timestamp 1666464484
transform 1 0 62944 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_558
timestamp 1666464484
transform 1 0 63840 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_560
timestamp 1666464484
transform 1 0 64064 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_575
timestamp 1666464484
transform 1 0 65744 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_591
timestamp 1666464484
transform 1 0 67536 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_599
timestamp 1666464484
transform 1 0 68432 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_605
timestamp 1666464484
transform 1 0 69104 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_669
timestamp 1666464484
transform 1 0 76272 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_673
timestamp 1666464484
transform 1 0 76720 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_676
timestamp 1666464484
transform 1 0 77056 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_740
timestamp 1666464484
transform 1 0 84224 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_744
timestamp 1666464484
transform 1 0 84672 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_747
timestamp 1666464484
transform 1 0 85008 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_755
timestamp 1666464484
transform 1 0 85904 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_759
timestamp 1666464484
transform 1 0 86352 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_761
timestamp 1666464484
transform 1 0 86576 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_764
timestamp 1666464484
transform 1 0 86912 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_772
timestamp 1666464484
transform 1 0 87808 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_804
timestamp 1666464484
transform 1 0 91392 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_812
timestamp 1666464484
transform 1 0 92288 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_818
timestamp 1666464484
transform 1 0 92960 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_882
timestamp 1666464484
transform 1 0 100128 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_886
timestamp 1666464484
transform 1 0 100576 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_889
timestamp 1666464484
transform 1 0 100912 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_953
timestamp 1666464484
transform 1 0 108080 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_957
timestamp 1666464484
transform 1 0 108528 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_960
timestamp 1666464484
transform 1 0 108864 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_968
timestamp 1666464484
transform 1 0 109760 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_972
timestamp 1666464484
transform 1 0 110208 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_976
timestamp 1666464484
transform 1 0 110656 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_1008
timestamp 1666464484
transform 1 0 114240 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1024
timestamp 1666464484
transform 1 0 116032 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1028
timestamp 1666464484
transform 1 0 116480 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_1031
timestamp 1666464484
transform 1 0 116816 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1095
timestamp 1666464484
transform 1 0 123984 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1099
timestamp 1666464484
transform 1 0 124432 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_1102
timestamp 1666464484
transform 1 0 124768 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1166
timestamp 1666464484
transform 1 0 131936 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1170
timestamp 1666464484
transform 1 0 132384 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_1173
timestamp 1666464484
transform 1 0 132720 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1237
timestamp 1666464484
transform 1 0 139888 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1241
timestamp 1666464484
transform 1 0 140336 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_1244
timestamp 1666464484
transform 1 0 140672 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1308
timestamp 1666464484
transform 1 0 147840 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1312
timestamp 1666464484
transform 1 0 148288 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_1315
timestamp 1666464484
transform 1 0 148624 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1379
timestamp 1666464484
transform 1 0 155792 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1383
timestamp 1666464484
transform 1 0 156240 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_1386
timestamp 1666464484
transform 1 0 156576 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1450
timestamp 1666464484
transform 1 0 163744 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1454
timestamp 1666464484
transform 1 0 164192 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_1457
timestamp 1666464484
transform 1 0 164528 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1521
timestamp 1666464484
transform 1 0 171696 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1525
timestamp 1666464484
transform 1 0 172144 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_1528
timestamp 1666464484
transform 1 0 172480 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_142_1560
timestamp 1666464484
transform 1 0 176064 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1576
timestamp 1666464484
transform 1 0 177856 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1580
timestamp 1666464484
transform 1 0 178304 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_2
timestamp 1666464484
transform 1 0 1568 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_18
timestamp 1666464484
transform 1 0 3360 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_32
timestamp 1666464484
transform 1 0 4928 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_36
timestamp 1666464484
transform 1 0 5376 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_44
timestamp 1666464484
transform 1 0 6272 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_46
timestamp 1666464484
transform 1 0 6496 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_49
timestamp 1666464484
transform 1 0 6832 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_57
timestamp 1666464484
transform 1 0 7728 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_61
timestamp 1666464484
transform 1 0 8176 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_69
timestamp 1666464484
transform 1 0 9072 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_73
timestamp 1666464484
transform 1 0 9520 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_81
timestamp 1666464484
transform 1 0 10416 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_85
timestamp 1666464484
transform 1 0 10864 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_89
timestamp 1666464484
transform 1 0 11312 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_97
timestamp 1666464484
transform 1 0 12208 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_113
timestamp 1666464484
transform 1 0 14000 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_129
timestamp 1666464484
transform 1 0 15792 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_133
timestamp 1666464484
transform 1 0 16240 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_141
timestamp 1666464484
transform 1 0 17136 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_144
timestamp 1666464484
transform 1 0 17472 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_159
timestamp 1666464484
transform 1 0 19152 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_167
timestamp 1666464484
transform 1 0 20048 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_171
timestamp 1666464484
transform 1 0 20496 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_173
timestamp 1666464484
transform 1 0 20720 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_176
timestamp 1666464484
transform 1 0 21056 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_184
timestamp 1666464484
transform 1 0 21952 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_200
timestamp 1666464484
transform 1 0 23744 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_208
timestamp 1666464484
transform 1 0 24640 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_212
timestamp 1666464484
transform 1 0 25088 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_215
timestamp 1666464484
transform 1 0 25424 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_218
timestamp 1666464484
transform 1 0 25760 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_226
timestamp 1666464484
transform 1 0 26656 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_260
timestamp 1666464484
transform 1 0 30464 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_268
timestamp 1666464484
transform 1 0 31360 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_272
timestamp 1666464484
transform 1 0 31808 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_280
timestamp 1666464484
transform 1 0 32704 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_286
timestamp 1666464484
transform 1 0 33376 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_294
timestamp 1666464484
transform 1 0 34272 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_296
timestamp 1666464484
transform 1 0 34496 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_299
timestamp 1666464484
transform 1 0 34832 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_307
timestamp 1666464484
transform 1 0 35728 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_323
timestamp 1666464484
transform 1 0 37520 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_339
timestamp 1666464484
transform 1 0 39312 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_341
timestamp 1666464484
transform 1 0 39536 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_344
timestamp 1666464484
transform 1 0 39872 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_352
timestamp 1666464484
transform 1 0 40768 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_354
timestamp 1666464484
transform 1 0 40992 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_357
timestamp 1666464484
transform 1 0 41328 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_372
timestamp 1666464484
transform 1 0 43008 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_380
timestamp 1666464484
transform 1 0 43904 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_386
timestamp 1666464484
transform 1 0 44576 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_394
timestamp 1666464484
transform 1 0 45472 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_410
timestamp 1666464484
transform 1 0 47264 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_418
timestamp 1666464484
transform 1 0 48160 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_422
timestamp 1666464484
transform 1 0 48608 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_425
timestamp 1666464484
transform 1 0 48944 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_428
timestamp 1666464484
transform 1 0 49280 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_436
timestamp 1666464484
transform 1 0 50176 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_470
timestamp 1666464484
transform 1 0 53984 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_478
timestamp 1666464484
transform 1 0 54880 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_482
timestamp 1666464484
transform 1 0 55328 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_490
timestamp 1666464484
transform 1 0 56224 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_494
timestamp 1666464484
transform 1 0 56672 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_496
timestamp 1666464484
transform 1 0 56896 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_499
timestamp 1666464484
transform 1 0 57232 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_509
timestamp 1666464484
transform 1 0 58352 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_517
timestamp 1666464484
transform 1 0 59248 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_533
timestamp 1666464484
transform 1 0 61040 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_549
timestamp 1666464484
transform 1 0 62832 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_551
timestamp 1666464484
transform 1 0 63056 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_554
timestamp 1666464484
transform 1 0 63392 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_562
timestamp 1666464484
transform 1 0 64288 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_566
timestamp 1666464484
transform 1 0 64736 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_570
timestamp 1666464484
transform 1 0 65184 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_586
timestamp 1666464484
transform 1 0 66976 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_596
timestamp 1666464484
transform 1 0 68096 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_604
timestamp 1666464484
transform 1 0 68992 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_638
timestamp 1666464484
transform 1 0 72800 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_641
timestamp 1666464484
transform 1 0 73136 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_648
timestamp 1666464484
transform 1 0 73920 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_664
timestamp 1666464484
transform 1 0 75712 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_672
timestamp 1666464484
transform 1 0 76608 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_676
timestamp 1666464484
transform 1 0 77056 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_680
timestamp 1666464484
transform 1 0 77504 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_688
timestamp 1666464484
transform 1 0 78400 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_692
timestamp 1666464484
transform 1 0 78848 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_708
timestamp 1666464484
transform 1 0 80640 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_712
timestamp 1666464484
transform 1 0 81088 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_716
timestamp 1666464484
transform 1 0 81536 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_719
timestamp 1666464484
transform 1 0 81872 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_727
timestamp 1666464484
transform 1 0 82768 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_743
timestamp 1666464484
transform 1 0 84560 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_759
timestamp 1666464484
transform 1 0 86352 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_763
timestamp 1666464484
transform 1 0 86800 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_765
timestamp 1666464484
transform 1 0 87024 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_780
timestamp 1666464484
transform 1 0 88704 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_783
timestamp 1666464484
transform 1 0 89040 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_799
timestamp 1666464484
transform 1 0 90832 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_803
timestamp 1666464484
transform 1 0 91280 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_806
timestamp 1666464484
transform 1 0 91616 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_814
timestamp 1666464484
transform 1 0 92512 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_822
timestamp 1666464484
transform 1 0 93408 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_826
timestamp 1666464484
transform 1 0 93856 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_841
timestamp 1666464484
transform 1 0 95536 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_845
timestamp 1666464484
transform 1 0 95984 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_851
timestamp 1666464484
transform 1 0 96656 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_854
timestamp 1666464484
transform 1 0 96992 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_861
timestamp 1666464484
transform 1 0 97776 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_877
timestamp 1666464484
transform 1 0 99568 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_885
timestamp 1666464484
transform 1 0 100464 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_887
timestamp 1666464484
transform 1 0 100688 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_890
timestamp 1666464484
transform 1 0 101024 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_898
timestamp 1666464484
transform 1 0 101920 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_902
timestamp 1666464484
transform 1 0 102368 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_918
timestamp 1666464484
transform 1 0 104160 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_922
timestamp 1666464484
transform 1 0 104608 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_925
timestamp 1666464484
transform 1 0 104944 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_931
timestamp 1666464484
transform 1 0 105616 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_939
timestamp 1666464484
transform 1 0 106512 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_947
timestamp 1666464484
transform 1 0 107408 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_951
timestamp 1666464484
transform 1 0 107856 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_967
timestamp 1666464484
transform 1 0 109648 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_971
timestamp 1666464484
transform 1 0 110096 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_975
timestamp 1666464484
transform 1 0 110544 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_982
timestamp 1666464484
transform 1 0 111328 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_990
timestamp 1666464484
transform 1 0 112224 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_996
timestamp 1666464484
transform 1 0 112896 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_999
timestamp 1666464484
transform 1 0 113232 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1007
timestamp 1666464484
transform 1 0 114128 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1011
timestamp 1666464484
transform 1 0 114576 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1013
timestamp 1666464484
transform 1 0 114800 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1016
timestamp 1666464484
transform 1 0 115136 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1024
timestamp 1666464484
transform 1 0 116032 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1032
timestamp 1666464484
transform 1 0 116928 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1035
timestamp 1666464484
transform 1 0 117264 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1051
timestamp 1666464484
transform 1 0 119056 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1059
timestamp 1666464484
transform 1 0 119952 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1061
timestamp 1666464484
transform 1 0 120176 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1064
timestamp 1666464484
transform 1 0 120512 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1067
timestamp 1666464484
transform 1 0 120848 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_1074
timestamp 1666464484
transform 1 0 121632 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1090
timestamp 1666464484
transform 1 0 123424 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1094
timestamp 1666464484
transform 1 0 123872 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1096
timestamp 1666464484
transform 1 0 124096 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1099
timestamp 1666464484
transform 1 0 124432 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1107
timestamp 1666464484
transform 1 0 125328 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1115
timestamp 1666464484
transform 1 0 126224 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1119
timestamp 1666464484
transform 1 0 126672 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1123
timestamp 1666464484
transform 1 0 127120 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1131
timestamp 1666464484
transform 1 0 128016 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1135
timestamp 1666464484
transform 1 0 128464 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1138
timestamp 1666464484
transform 1 0 128800 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1141
timestamp 1666464484
transform 1 0 129136 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1149
timestamp 1666464484
transform 1 0 130032 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1157
timestamp 1666464484
transform 1 0 130928 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1161
timestamp 1666464484
transform 1 0 131376 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1177
timestamp 1666464484
transform 1 0 133168 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1181
timestamp 1666464484
transform 1 0 133616 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1184
timestamp 1666464484
transform 1 0 133952 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1192
timestamp 1666464484
transform 1 0 134848 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1200
timestamp 1666464484
transform 1 0 135744 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1204
timestamp 1666464484
transform 1 0 136192 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1206
timestamp 1666464484
transform 1 0 136416 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1209
timestamp 1666464484
transform 1 0 136752 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1212
timestamp 1666464484
transform 1 0 137088 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1220
timestamp 1666464484
transform 1 0 137984 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1226
timestamp 1666464484
transform 1 0 138656 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1234
timestamp 1666464484
transform 1 0 139552 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1242
timestamp 1666464484
transform 1 0 140448 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1245
timestamp 1666464484
transform 1 0 140784 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1261
timestamp 1666464484
transform 1 0 142576 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1265
timestamp 1666464484
transform 1 0 143024 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1268
timestamp 1666464484
transform 1 0 143360 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1276
timestamp 1666464484
transform 1 0 144256 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_1280
timestamp 1666464484
transform 1 0 144704 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1296
timestamp 1666464484
transform 1 0 146496 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1304
timestamp 1666464484
transform 1 0 147392 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1310
timestamp 1666464484
transform 1 0 148064 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1318
timestamp 1666464484
transform 1 0 148960 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1326
timestamp 1666464484
transform 1 0 149856 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1330
timestamp 1666464484
transform 1 0 150304 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1333
timestamp 1666464484
transform 1 0 150640 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1341
timestamp 1666464484
transform 1 0 151536 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1345
timestamp 1666464484
transform 1 0 151984 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1348
timestamp 1666464484
transform 1 0 152320 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1351
timestamp 1666464484
transform 1 0 152656 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1353
timestamp 1666464484
transform 1 0 152880 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1360
timestamp 1666464484
transform 1 0 153664 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1368
timestamp 1666464484
transform 1 0 154560 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1372
timestamp 1666464484
transform 1 0 155008 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1377
timestamp 1666464484
transform 1 0 155568 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1385
timestamp 1666464484
transform 1 0 156464 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1389
timestamp 1666464484
transform 1 0 156912 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1391
timestamp 1666464484
transform 1 0 157136 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1394
timestamp 1666464484
transform 1 0 157472 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_143_1402
timestamp 1666464484
transform 1 0 158368 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1418
timestamp 1666464484
transform 1 0 160160 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1422
timestamp 1666464484
transform 1 0 160608 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1430
timestamp 1666464484
transform 1 0 161504 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1436
timestamp 1666464484
transform 1 0 162176 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_1444
timestamp 1666464484
transform 1 0 163072 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1478
timestamp 1666464484
transform 1 0 166880 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1486
timestamp 1666464484
transform 1 0 167776 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1490
timestamp 1666464484
transform 1 0 168224 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1493
timestamp 1666464484
transform 1 0 168560 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1501
timestamp 1666464484
transform 1 0 169456 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1505
timestamp 1666464484
transform 1 0 169904 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1508
timestamp 1666464484
transform 1 0 170240 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_1516
timestamp 1666464484
transform 1 0 171136 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1548
timestamp 1666464484
transform 1 0 174720 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1556
timestamp 1666464484
transform 1 0 175616 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_1560
timestamp 1666464484
transform 1 0 176064 0 -1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1564
timestamp 1666464484
transform 1 0 176512 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1572
timestamp 1666464484
transform 1 0 177408 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1580
timestamp 1666464484
transform 1 0 178304 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_2
timestamp 1666464484
transform 1 0 1568 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_10
timestamp 1666464484
transform 1 0 2464 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_14
timestamp 1666464484
transform 1 0 2912 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_29
timestamp 1666464484
transform 1 0 4592 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_33
timestamp 1666464484
transform 1 0 5040 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_37
timestamp 1666464484
transform 1 0 5488 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_52
timestamp 1666464484
transform 1 0 7168 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_54
timestamp 1666464484
transform 1 0 7392 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_69
timestamp 1666464484
transform 1 0 9072 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_72
timestamp 1666464484
transform 1 0 9408 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_87
timestamp 1666464484
transform 1 0 11088 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_91
timestamp 1666464484
transform 1 0 11536 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_99
timestamp 1666464484
transform 1 0 12432 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_103
timestamp 1666464484
transform 1 0 12880 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_107
timestamp 1666464484
transform 1 0 13328 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_111
timestamp 1666464484
transform 1 0 13776 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_127
timestamp 1666464484
transform 1 0 15568 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_131
timestamp 1666464484
transform 1 0 16016 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_139
timestamp 1666464484
transform 1 0 16912 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_142
timestamp 1666464484
transform 1 0 17248 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_150
timestamp 1666464484
transform 1 0 18144 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_154
timestamp 1666464484
transform 1 0 18592 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_169
timestamp 1666464484
transform 1 0 20272 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_173
timestamp 1666464484
transform 1 0 20720 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_177
timestamp 1666464484
transform 1 0 21168 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_193
timestamp 1666464484
transform 1 0 22960 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_209
timestamp 1666464484
transform 1 0 24752 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_212
timestamp 1666464484
transform 1 0 25088 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_215
timestamp 1666464484
transform 1 0 25424 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_223
timestamp 1666464484
transform 1 0 26320 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_239
timestamp 1666464484
transform 1 0 28112 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_243
timestamp 1666464484
transform 1 0 28560 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_247
timestamp 1666464484
transform 1 0 29008 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_262
timestamp 1666464484
transform 1 0 30688 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_264
timestamp 1666464484
transform 1 0 30912 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_279
timestamp 1666464484
transform 1 0 32592 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_282
timestamp 1666464484
transform 1 0 32928 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_297
timestamp 1666464484
transform 1 0 34608 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_301
timestamp 1666464484
transform 1 0 35056 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_309
timestamp 1666464484
transform 1 0 35952 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_313
timestamp 1666464484
transform 1 0 36400 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_317
timestamp 1666464484
transform 1 0 36848 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_321
timestamp 1666464484
transform 1 0 37296 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_337
timestamp 1666464484
transform 1 0 39088 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_341
timestamp 1666464484
transform 1 0 39536 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_349
timestamp 1666464484
transform 1 0 40432 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_352
timestamp 1666464484
transform 1 0 40768 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_360
timestamp 1666464484
transform 1 0 41664 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_364
timestamp 1666464484
transform 1 0 42112 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_379
timestamp 1666464484
transform 1 0 43792 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_383
timestamp 1666464484
transform 1 0 44240 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_387
timestamp 1666464484
transform 1 0 44688 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_403
timestamp 1666464484
transform 1 0 46480 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_419
timestamp 1666464484
transform 1 0 48272 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_422
timestamp 1666464484
transform 1 0 48608 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_425
timestamp 1666464484
transform 1 0 48944 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_433
timestamp 1666464484
transform 1 0 49840 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_449
timestamp 1666464484
transform 1 0 51632 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_453
timestamp 1666464484
transform 1 0 52080 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_457
timestamp 1666464484
transform 1 0 52528 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_472
timestamp 1666464484
transform 1 0 54208 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_474
timestamp 1666464484
transform 1 0 54432 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_489
timestamp 1666464484
transform 1 0 56112 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_492
timestamp 1666464484
transform 1 0 56448 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_507
timestamp 1666464484
transform 1 0 58128 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_511
timestamp 1666464484
transform 1 0 58576 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_519
timestamp 1666464484
transform 1 0 59472 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_523
timestamp 1666464484
transform 1 0 59920 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_527
timestamp 1666464484
transform 1 0 60368 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_531
timestamp 1666464484
transform 1 0 60816 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_547
timestamp 1666464484
transform 1 0 62608 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_551
timestamp 1666464484
transform 1 0 63056 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_559
timestamp 1666464484
transform 1 0 63952 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_562
timestamp 1666464484
transform 1 0 64288 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_570
timestamp 1666464484
transform 1 0 65184 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_574
timestamp 1666464484
transform 1 0 65632 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_589
timestamp 1666464484
transform 1 0 67312 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_593
timestamp 1666464484
transform 1 0 67760 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_597
timestamp 1666464484
transform 1 0 68208 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_613
timestamp 1666464484
transform 1 0 70000 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_629
timestamp 1666464484
transform 1 0 71792 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_632
timestamp 1666464484
transform 1 0 72128 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_635
timestamp 1666464484
transform 1 0 72464 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_643
timestamp 1666464484
transform 1 0 73360 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_659
timestamp 1666464484
transform 1 0 75152 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_663
timestamp 1666464484
transform 1 0 75600 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_667
timestamp 1666464484
transform 1 0 76048 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_682
timestamp 1666464484
transform 1 0 77728 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_684
timestamp 1666464484
transform 1 0 77952 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_699
timestamp 1666464484
transform 1 0 79632 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_702
timestamp 1666464484
transform 1 0 79968 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_717
timestamp 1666464484
transform 1 0 81648 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_721
timestamp 1666464484
transform 1 0 82096 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_729
timestamp 1666464484
transform 1 0 82992 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_733
timestamp 1666464484
transform 1 0 83440 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_737
timestamp 1666464484
transform 1 0 83888 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_741
timestamp 1666464484
transform 1 0 84336 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_757
timestamp 1666464484
transform 1 0 86128 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_761
timestamp 1666464484
transform 1 0 86576 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_769
timestamp 1666464484
transform 1 0 87472 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_772
timestamp 1666464484
transform 1 0 87808 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_780
timestamp 1666464484
transform 1 0 88704 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_784
timestamp 1666464484
transform 1 0 89152 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_799
timestamp 1666464484
transform 1 0 90832 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_803
timestamp 1666464484
transform 1 0 91280 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_807
timestamp 1666464484
transform 1 0 91728 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_811
timestamp 1666464484
transform 1 0 92176 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_827
timestamp 1666464484
transform 1 0 93968 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_835
timestamp 1666464484
transform 1 0 94864 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_839
timestamp 1666464484
transform 1 0 95312 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_842
timestamp 1666464484
transform 1 0 95648 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_850
timestamp 1666464484
transform 1 0 96544 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_854
timestamp 1666464484
transform 1 0 96992 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_869
timestamp 1666464484
transform 1 0 98672 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_873
timestamp 1666464484
transform 1 0 99120 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_877
timestamp 1666464484
transform 1 0 99568 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_892
timestamp 1666464484
transform 1 0 101248 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_894
timestamp 1666464484
transform 1 0 101472 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_909
timestamp 1666464484
transform 1 0 103152 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_912
timestamp 1666464484
transform 1 0 103488 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_927
timestamp 1666464484
transform 1 0 105168 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_931
timestamp 1666464484
transform 1 0 105616 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_939
timestamp 1666464484
transform 1 0 106512 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_943
timestamp 1666464484
transform 1 0 106960 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_947
timestamp 1666464484
transform 1 0 107408 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_962
timestamp 1666464484
transform 1 0 109088 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_978
timestamp 1666464484
transform 1 0 110880 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_982
timestamp 1666464484
transform 1 0 111328 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_997
timestamp 1666464484
transform 1 0 113008 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1013
timestamp 1666464484
transform 1 0 114800 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1017
timestamp 1666464484
transform 1 0 115248 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1021
timestamp 1666464484
transform 1 0 115696 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1037
timestamp 1666464484
transform 1 0 117488 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1045
timestamp 1666464484
transform 1 0 118384 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1049
timestamp 1666464484
transform 1 0 118832 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1052
timestamp 1666464484
transform 1 0 119168 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1060
timestamp 1666464484
transform 1 0 120064 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1064
timestamp 1666464484
transform 1 0 120512 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1079
timestamp 1666464484
transform 1 0 122192 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1081
timestamp 1666464484
transform 1 0 122416 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1084
timestamp 1666464484
transform 1 0 122752 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1087
timestamp 1666464484
transform 1 0 123088 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1102
timestamp 1666464484
transform 1 0 124768 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1104
timestamp 1666464484
transform 1 0 124992 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1119
timestamp 1666464484
transform 1 0 126672 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1122
timestamp 1666464484
transform 1 0 127008 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_1137
timestamp 1666464484
transform 1 0 128688 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1153
timestamp 1666464484
transform 1 0 130480 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1157
timestamp 1666464484
transform 1 0 130928 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_1172
timestamp 1666464484
transform 1 0 132608 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1188
timestamp 1666464484
transform 1 0 134400 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1192
timestamp 1666464484
transform 1 0 134848 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1207
timestamp 1666464484
transform 1 0 136528 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1223
timestamp 1666464484
transform 1 0 138320 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1227
timestamp 1666464484
transform 1 0 138768 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1231
timestamp 1666464484
transform 1 0 139216 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1247
timestamp 1666464484
transform 1 0 141008 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1255
timestamp 1666464484
transform 1 0 141904 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1259
timestamp 1666464484
transform 1 0 142352 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1262
timestamp 1666464484
transform 1 0 142688 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1270
timestamp 1666464484
transform 1 0 143584 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1274
timestamp 1666464484
transform 1 0 144032 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1289
timestamp 1666464484
transform 1 0 145712 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1291
timestamp 1666464484
transform 1 0 145936 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1294
timestamp 1666464484
transform 1 0 146272 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1297
timestamp 1666464484
transform 1 0 146608 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1312
timestamp 1666464484
transform 1 0 148288 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1314
timestamp 1666464484
transform 1 0 148512 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1329
timestamp 1666464484
transform 1 0 150192 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1332
timestamp 1666464484
transform 1 0 150528 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_1347
timestamp 1666464484
transform 1 0 152208 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1363
timestamp 1666464484
transform 1 0 154000 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1367
timestamp 1666464484
transform 1 0 154448 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_1382
timestamp 1666464484
transform 1 0 156128 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1398
timestamp 1666464484
transform 1 0 157920 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1402
timestamp 1666464484
transform 1 0 158368 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1417
timestamp 1666464484
transform 1 0 160048 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1423
timestamp 1666464484
transform 1 0 160720 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1431
timestamp 1666464484
transform 1 0 161616 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1437
timestamp 1666464484
transform 1 0 162288 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1441
timestamp 1666464484
transform 1 0 162736 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1457
timestamp 1666464484
transform 1 0 164528 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1463
timestamp 1666464484
transform 1 0 165200 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1467
timestamp 1666464484
transform 1 0 165648 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1469
timestamp 1666464484
transform 1 0 165872 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1472
timestamp 1666464484
transform 1 0 166208 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1480
timestamp 1666464484
transform 1 0 167104 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1484
timestamp 1666464484
transform 1 0 167552 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1499
timestamp 1666464484
transform 1 0 169232 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1503
timestamp 1666464484
transform 1 0 169680 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1507
timestamp 1666464484
transform 1 0 170128 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1512
timestamp 1666464484
transform 1 0 170688 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1520
timestamp 1666464484
transform 1 0 171584 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1524
timestamp 1666464484
transform 1 0 172032 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1539
timestamp 1666464484
transform 1 0 173712 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1542
timestamp 1666464484
transform 1 0 174048 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_144_1547
timestamp 1666464484
transform 1 0 174608 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1563
timestamp 1666464484
transform 1 0 176400 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1567
timestamp 1666464484
transform 1 0 176848 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_144_1573
timestamp 1666464484
transform 1 0 177520 0 1 116032
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1577
timestamp 1666464484
transform 1 0 177968 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 178640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 178640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 178640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 178640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 178640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 178640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 178640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 178640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 178640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 178640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 178640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1666464484
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1666464484
transform -1 0 178640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1666464484
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1666464484
transform -1 0 178640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1666464484
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1666464484
transform -1 0 178640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1666464484
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1666464484
transform -1 0 178640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1666464484
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1666464484
transform -1 0 178640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1666464484
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1666464484
transform -1 0 178640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1666464484
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1666464484
transform -1 0 178640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1666464484
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1666464484
transform -1 0 178640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1666464484
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1666464484
transform -1 0 178640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1666464484
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1666464484
transform -1 0 178640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1666464484
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1666464484
transform -1 0 178640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1666464484
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1666464484
transform -1 0 178640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1666464484
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1666464484
transform -1 0 178640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1666464484
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1666464484
transform -1 0 178640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1666464484
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1666464484
transform -1 0 178640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1666464484
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1666464484
transform -1 0 178640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1666464484
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1666464484
transform -1 0 178640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1666464484
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1666464484
transform -1 0 178640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1666464484
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1666464484
transform -1 0 178640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1666464484
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1666464484
transform -1 0 178640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1666464484
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1666464484
transform -1 0 178640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1666464484
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1666464484
transform -1 0 178640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1666464484
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1666464484
transform -1 0 178640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1666464484
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1666464484
transform -1 0 178640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1666464484
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1666464484
transform -1 0 178640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1666464484
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1666464484
transform -1 0 178640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1666464484
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1666464484
transform -1 0 178640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1666464484
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1666464484
transform -1 0 178640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1666464484
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1666464484
transform -1 0 178640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1666464484
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1666464484
transform -1 0 178640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1666464484
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1666464484
transform -1 0 178640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1666464484
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1666464484
transform -1 0 178640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1666464484
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1666464484
transform -1 0 178640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1666464484
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1666464484
transform -1 0 178640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1666464484
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1666464484
transform -1 0 178640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1666464484
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1666464484
transform -1 0 178640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1666464484
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1666464484
transform -1 0 178640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1666464484
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1666464484
transform -1 0 178640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1666464484
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1666464484
transform -1 0 178640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1666464484
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1666464484
transform -1 0 178640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1666464484
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1666464484
transform -1 0 178640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1666464484
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1666464484
transform -1 0 178640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1666464484
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1666464484
transform -1 0 178640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1666464484
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1666464484
transform -1 0 178640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1666464484
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1666464484
transform -1 0 178640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1666464484
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1666464484
transform -1 0 178640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1666464484
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1666464484
transform -1 0 178640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1666464484
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1666464484
transform -1 0 178640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1666464484
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1666464484
transform -1 0 178640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1666464484
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1666464484
transform -1 0 178640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1666464484
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1666464484
transform -1 0 178640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1666464484
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1666464484
transform -1 0 178640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1666464484
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1666464484
transform -1 0 178640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1666464484
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1666464484
transform -1 0 178640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1666464484
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1666464484
transform -1 0 178640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1666464484
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1666464484
transform -1 0 178640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1666464484
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1666464484
transform -1 0 178640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1666464484
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1666464484
transform -1 0 178640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1666464484
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1666464484
transform -1 0 178640 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1666464484
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1666464484
transform -1 0 178640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1666464484
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1666464484
transform -1 0 178640 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1666464484
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1666464484
transform -1 0 178640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1666464484
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1666464484
transform -1 0 178640 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1666464484
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1666464484
transform -1 0 178640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1666464484
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1666464484
transform -1 0 178640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1666464484
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1666464484
transform -1 0 178640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1666464484
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1666464484
transform -1 0 178640 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1666464484
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1666464484
transform -1 0 178640 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1666464484
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1666464484
transform -1 0 178640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1666464484
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1666464484
transform -1 0 178640 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1666464484
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1666464484
transform -1 0 178640 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1666464484
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1666464484
transform -1 0 178640 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1666464484
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1666464484
transform -1 0 178640 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1666464484
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1666464484
transform -1 0 178640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1666464484
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1666464484
transform -1 0 178640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1666464484
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1666464484
transform -1 0 178640 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1666464484
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1666464484
transform -1 0 178640 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1666464484
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1666464484
transform -1 0 178640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1666464484
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1666464484
transform -1 0 178640 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1666464484
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1666464484
transform -1 0 178640 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1666464484
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1666464484
transform -1 0 178640 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1666464484
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1666464484
transform -1 0 178640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1666464484
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1666464484
transform -1 0 178640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_188
timestamp 1666464484
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_189
timestamp 1666464484
transform -1 0 178640 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_190
timestamp 1666464484
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_191
timestamp 1666464484
transform -1 0 178640 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_192
timestamp 1666464484
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_193
timestamp 1666464484
transform -1 0 178640 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_194
timestamp 1666464484
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_195
timestamp 1666464484
transform -1 0 178640 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_196
timestamp 1666464484
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_197
timestamp 1666464484
transform -1 0 178640 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_198
timestamp 1666464484
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_199
timestamp 1666464484
transform -1 0 178640 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_200
timestamp 1666464484
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_201
timestamp 1666464484
transform -1 0 178640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_202
timestamp 1666464484
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_203
timestamp 1666464484
transform -1 0 178640 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_204
timestamp 1666464484
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_205
timestamp 1666464484
transform -1 0 178640 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_206
timestamp 1666464484
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_207
timestamp 1666464484
transform -1 0 178640 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_208
timestamp 1666464484
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_209
timestamp 1666464484
transform -1 0 178640 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_210
timestamp 1666464484
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_211
timestamp 1666464484
transform -1 0 178640 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_212
timestamp 1666464484
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_213
timestamp 1666464484
transform -1 0 178640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_214
timestamp 1666464484
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_215
timestamp 1666464484
transform -1 0 178640 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_216
timestamp 1666464484
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_217
timestamp 1666464484
transform -1 0 178640 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_218
timestamp 1666464484
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_219
timestamp 1666464484
transform -1 0 178640 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_220
timestamp 1666464484
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_221
timestamp 1666464484
transform -1 0 178640 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_222
timestamp 1666464484
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_223
timestamp 1666464484
transform -1 0 178640 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_224
timestamp 1666464484
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_225
timestamp 1666464484
transform -1 0 178640 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_226
timestamp 1666464484
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_227
timestamp 1666464484
transform -1 0 178640 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_228
timestamp 1666464484
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_229
timestamp 1666464484
transform -1 0 178640 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_230
timestamp 1666464484
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_231
timestamp 1666464484
transform -1 0 178640 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_232
timestamp 1666464484
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_233
timestamp 1666464484
transform -1 0 178640 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_234
timestamp 1666464484
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_235
timestamp 1666464484
transform -1 0 178640 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_236
timestamp 1666464484
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_237
timestamp 1666464484
transform -1 0 178640 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_238
timestamp 1666464484
transform 1 0 1344 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_239
timestamp 1666464484
transform -1 0 178640 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_240
timestamp 1666464484
transform 1 0 1344 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_241
timestamp 1666464484
transform -1 0 178640 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_242
timestamp 1666464484
transform 1 0 1344 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_243
timestamp 1666464484
transform -1 0 178640 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_244
timestamp 1666464484
transform 1 0 1344 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_245
timestamp 1666464484
transform -1 0 178640 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_246
timestamp 1666464484
transform 1 0 1344 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_247
timestamp 1666464484
transform -1 0 178640 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_248
timestamp 1666464484
transform 1 0 1344 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_249
timestamp 1666464484
transform -1 0 178640 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_250
timestamp 1666464484
transform 1 0 1344 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_251
timestamp 1666464484
transform -1 0 178640 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_252
timestamp 1666464484
transform 1 0 1344 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_253
timestamp 1666464484
transform -1 0 178640 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_254
timestamp 1666464484
transform 1 0 1344 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_255
timestamp 1666464484
transform -1 0 178640 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_256
timestamp 1666464484
transform 1 0 1344 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_257
timestamp 1666464484
transform -1 0 178640 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_258
timestamp 1666464484
transform 1 0 1344 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_259
timestamp 1666464484
transform -1 0 178640 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_260
timestamp 1666464484
transform 1 0 1344 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_261
timestamp 1666464484
transform -1 0 178640 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_262
timestamp 1666464484
transform 1 0 1344 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_263
timestamp 1666464484
transform -1 0 178640 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_264
timestamp 1666464484
transform 1 0 1344 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_265
timestamp 1666464484
transform -1 0 178640 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_266
timestamp 1666464484
transform 1 0 1344 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_267
timestamp 1666464484
transform -1 0 178640 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_268
timestamp 1666464484
transform 1 0 1344 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_269
timestamp 1666464484
transform -1 0 178640 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_270
timestamp 1666464484
transform 1 0 1344 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_271
timestamp 1666464484
transform -1 0 178640 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_272
timestamp 1666464484
transform 1 0 1344 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_273
timestamp 1666464484
transform -1 0 178640 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_274
timestamp 1666464484
transform 1 0 1344 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_275
timestamp 1666464484
transform -1 0 178640 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_276
timestamp 1666464484
transform 1 0 1344 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_277
timestamp 1666464484
transform -1 0 178640 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_278
timestamp 1666464484
transform 1 0 1344 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_279
timestamp 1666464484
transform -1 0 178640 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_280
timestamp 1666464484
transform 1 0 1344 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_281
timestamp 1666464484
transform -1 0 178640 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_282
timestamp 1666464484
transform 1 0 1344 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_283
timestamp 1666464484
transform -1 0 178640 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_284
timestamp 1666464484
transform 1 0 1344 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_285
timestamp 1666464484
transform -1 0 178640 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_286
timestamp 1666464484
transform 1 0 1344 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_287
timestamp 1666464484
transform -1 0 178640 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_288
timestamp 1666464484
transform 1 0 1344 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_289
timestamp 1666464484
transform -1 0 178640 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1666464484
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1666464484
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1666464484
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1666464484
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1666464484
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1666464484
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1666464484
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1666464484
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1666464484
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1666464484
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1666464484
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1666464484
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1666464484
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1666464484
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1666464484
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1666464484
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1666464484
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1666464484
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1666464484
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1666464484
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1666464484
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1666464484
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1666464484
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1666464484
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1666464484
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1666464484
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1666464484
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1666464484
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1666464484
transform 1 0 118944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1666464484
transform 1 0 122864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1666464484
transform 1 0 126784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1666464484
transform 1 0 130704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1666464484
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1666464484
transform 1 0 138544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1666464484
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1666464484
transform 1 0 146384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1666464484
transform 1 0 150304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1666464484
transform 1 0 154224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1666464484
transform 1 0 158144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1666464484
transform 1 0 162064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1666464484
transform 1 0 165984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1666464484
transform 1 0 169904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1666464484
transform 1 0 173824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1666464484
transform 1 0 177744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1666464484
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1666464484
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1666464484
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1666464484
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1666464484
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1666464484
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1666464484
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1666464484
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1666464484
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1666464484
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1666464484
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1666464484
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1666464484
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1666464484
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1666464484
transform 1 0 120624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1666464484
transform 1 0 128576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1666464484
transform 1 0 136528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1666464484
transform 1 0 144480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1666464484
transform 1 0 152432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1666464484
transform 1 0 160384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1666464484
transform 1 0 168336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1666464484
transform 1 0 176288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1666464484
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1666464484
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1666464484
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1666464484
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1666464484
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1666464484
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1666464484
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1666464484
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1666464484
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1666464484
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1666464484
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1666464484
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1666464484
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1666464484
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1666464484
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1666464484
transform 1 0 124544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1666464484
transform 1 0 132496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1666464484
transform 1 0 140448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1666464484
transform 1 0 148400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1666464484
transform 1 0 156352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1666464484
transform 1 0 164304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1666464484
transform 1 0 172256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1666464484
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1666464484
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1666464484
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1666464484
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1666464484
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1666464484
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1666464484
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1666464484
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1666464484
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1666464484
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1666464484
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1666464484
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1666464484
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1666464484
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1666464484
transform 1 0 120624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1666464484
transform 1 0 128576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1666464484
transform 1 0 136528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1666464484
transform 1 0 144480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1666464484
transform 1 0 152432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1666464484
transform 1 0 160384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1666464484
transform 1 0 168336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1666464484
transform 1 0 176288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1666464484
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1666464484
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1666464484
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1666464484
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1666464484
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1666464484
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1666464484
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1666464484
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1666464484
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1666464484
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1666464484
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1666464484
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1666464484
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1666464484
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1666464484
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1666464484
transform 1 0 124544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1666464484
transform 1 0 132496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1666464484
transform 1 0 140448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1666464484
transform 1 0 148400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1666464484
transform 1 0 156352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1666464484
transform 1 0 164304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1666464484
transform 1 0 172256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1666464484
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1666464484
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1666464484
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1666464484
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1666464484
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1666464484
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1666464484
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1666464484
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1666464484
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1666464484
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1666464484
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1666464484
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1666464484
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1666464484
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1666464484
transform 1 0 120624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1666464484
transform 1 0 128576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1666464484
transform 1 0 136528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1666464484
transform 1 0 144480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1666464484
transform 1 0 152432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1666464484
transform 1 0 160384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1666464484
transform 1 0 168336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1666464484
transform 1 0 176288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1666464484
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1666464484
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1666464484
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1666464484
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1666464484
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1666464484
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1666464484
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1666464484
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1666464484
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1666464484
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1666464484
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1666464484
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1666464484
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1666464484
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1666464484
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1666464484
transform 1 0 124544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1666464484
transform 1 0 132496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1666464484
transform 1 0 140448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1666464484
transform 1 0 148400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1666464484
transform 1 0 156352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1666464484
transform 1 0 164304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1666464484
transform 1 0 172256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1666464484
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1666464484
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1666464484
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1666464484
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1666464484
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1666464484
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1666464484
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1666464484
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1666464484
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1666464484
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1666464484
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1666464484
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1666464484
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1666464484
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1666464484
transform 1 0 120624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1666464484
transform 1 0 128576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1666464484
transform 1 0 136528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1666464484
transform 1 0 144480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1666464484
transform 1 0 152432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1666464484
transform 1 0 160384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1666464484
transform 1 0 168336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1666464484
transform 1 0 176288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1666464484
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1666464484
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1666464484
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1666464484
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1666464484
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1666464484
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1666464484
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1666464484
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1666464484
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1666464484
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1666464484
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1666464484
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1666464484
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1666464484
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1666464484
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1666464484
transform 1 0 124544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1666464484
transform 1 0 132496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1666464484
transform 1 0 140448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1666464484
transform 1 0 148400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1666464484
transform 1 0 156352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1666464484
transform 1 0 164304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1666464484
transform 1 0 172256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1666464484
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1666464484
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1666464484
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1666464484
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1666464484
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1666464484
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1666464484
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1666464484
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1666464484
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1666464484
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1666464484
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1666464484
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1666464484
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1666464484
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1666464484
transform 1 0 120624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1666464484
transform 1 0 128576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1666464484
transform 1 0 136528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1666464484
transform 1 0 144480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1666464484
transform 1 0 152432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1666464484
transform 1 0 160384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1666464484
transform 1 0 168336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1666464484
transform 1 0 176288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1666464484
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1666464484
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1666464484
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1666464484
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1666464484
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1666464484
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1666464484
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1666464484
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1666464484
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1666464484
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1666464484
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1666464484
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1666464484
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1666464484
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1666464484
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1666464484
transform 1 0 124544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1666464484
transform 1 0 132496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1666464484
transform 1 0 140448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1666464484
transform 1 0 148400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1666464484
transform 1 0 156352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1666464484
transform 1 0 164304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1666464484
transform 1 0 172256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1666464484
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1666464484
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1666464484
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1666464484
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1666464484
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1666464484
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1666464484
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1666464484
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1666464484
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1666464484
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1666464484
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1666464484
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1666464484
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1666464484
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1666464484
transform 1 0 120624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1666464484
transform 1 0 128576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1666464484
transform 1 0 136528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1666464484
transform 1 0 144480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1666464484
transform 1 0 152432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1666464484
transform 1 0 160384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1666464484
transform 1 0 168336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1666464484
transform 1 0 176288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1666464484
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1666464484
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1666464484
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1666464484
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1666464484
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1666464484
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1666464484
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1666464484
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1666464484
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1666464484
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1666464484
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1666464484
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1666464484
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1666464484
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1666464484
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1666464484
transform 1 0 124544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1666464484
transform 1 0 132496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1666464484
transform 1 0 140448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1666464484
transform 1 0 148400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1666464484
transform 1 0 156352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1666464484
transform 1 0 164304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1666464484
transform 1 0 172256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1666464484
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1666464484
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1666464484
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1666464484
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1666464484
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1666464484
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1666464484
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1666464484
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1666464484
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1666464484
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1666464484
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1666464484
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1666464484
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1666464484
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1666464484
transform 1 0 120624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1666464484
transform 1 0 128576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1666464484
transform 1 0 136528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1666464484
transform 1 0 144480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1666464484
transform 1 0 152432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1666464484
transform 1 0 160384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1666464484
transform 1 0 168336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1666464484
transform 1 0 176288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1666464484
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1666464484
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1666464484
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1666464484
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1666464484
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1666464484
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1666464484
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1666464484
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1666464484
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1666464484
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1666464484
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1666464484
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1666464484
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1666464484
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1666464484
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1666464484
transform 1 0 124544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1666464484
transform 1 0 132496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1666464484
transform 1 0 140448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1666464484
transform 1 0 148400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1666464484
transform 1 0 156352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1666464484
transform 1 0 164304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1666464484
transform 1 0 172256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1666464484
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1666464484
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1666464484
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1666464484
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1666464484
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1666464484
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1666464484
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1666464484
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1666464484
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1666464484
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1666464484
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1666464484
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1666464484
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1666464484
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1666464484
transform 1 0 120624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1666464484
transform 1 0 128576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1666464484
transform 1 0 136528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1666464484
transform 1 0 144480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1666464484
transform 1 0 152432 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1666464484
transform 1 0 160384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1666464484
transform 1 0 168336 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1666464484
transform 1 0 176288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1666464484
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1666464484
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1666464484
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1666464484
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1666464484
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1666464484
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1666464484
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1666464484
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1666464484
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1666464484
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1666464484
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1666464484
transform 1 0 92736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1666464484
transform 1 0 100688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1666464484
transform 1 0 108640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1666464484
transform 1 0 116592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1666464484
transform 1 0 124544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1666464484
transform 1 0 132496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1666464484
transform 1 0 140448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1666464484
transform 1 0 148400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1666464484
transform 1 0 156352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1666464484
transform 1 0 164304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1666464484
transform 1 0 172256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1666464484
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1666464484
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1666464484
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1666464484
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1666464484
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1666464484
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1666464484
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1666464484
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1666464484
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1666464484
transform 1 0 80864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1666464484
transform 1 0 88816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1666464484
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1666464484
transform 1 0 104720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1666464484
transform 1 0 112672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1666464484
transform 1 0 120624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1666464484
transform 1 0 128576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1666464484
transform 1 0 136528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1666464484
transform 1 0 144480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1666464484
transform 1 0 152432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1666464484
transform 1 0 160384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1666464484
transform 1 0 168336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1666464484
transform 1 0 176288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1666464484
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1666464484
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1666464484
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1666464484
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1666464484
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1666464484
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1666464484
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1666464484
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1666464484
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1666464484
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1666464484
transform 1 0 84784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1666464484
transform 1 0 92736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1666464484
transform 1 0 100688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1666464484
transform 1 0 108640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1666464484
transform 1 0 116592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1666464484
transform 1 0 124544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1666464484
transform 1 0 132496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1666464484
transform 1 0 140448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1666464484
transform 1 0 148400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1666464484
transform 1 0 156352 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1666464484
transform 1 0 164304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1666464484
transform 1 0 172256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1666464484
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1666464484
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1666464484
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1666464484
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1666464484
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1666464484
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1666464484
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1666464484
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1666464484
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1666464484
transform 1 0 80864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1666464484
transform 1 0 88816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1666464484
transform 1 0 96768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1666464484
transform 1 0 104720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1666464484
transform 1 0 112672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1666464484
transform 1 0 120624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1666464484
transform 1 0 128576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1666464484
transform 1 0 136528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1666464484
transform 1 0 144480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1666464484
transform 1 0 152432 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1666464484
transform 1 0 160384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1666464484
transform 1 0 168336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1666464484
transform 1 0 176288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1666464484
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1666464484
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1666464484
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1666464484
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1666464484
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1666464484
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1666464484
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1666464484
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1666464484
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1666464484
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1666464484
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1666464484
transform 1 0 92736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1666464484
transform 1 0 100688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1666464484
transform 1 0 108640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1666464484
transform 1 0 116592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1666464484
transform 1 0 124544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1666464484
transform 1 0 132496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1666464484
transform 1 0 140448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1666464484
transform 1 0 148400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1666464484
transform 1 0 156352 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1666464484
transform 1 0 164304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1666464484
transform 1 0 172256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1666464484
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1666464484
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1666464484
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1666464484
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1666464484
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1666464484
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1666464484
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1666464484
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1666464484
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1666464484
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1666464484
transform 1 0 88816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1666464484
transform 1 0 96768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1666464484
transform 1 0 104720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1666464484
transform 1 0 112672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1666464484
transform 1 0 120624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1666464484
transform 1 0 128576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1666464484
transform 1 0 136528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1666464484
transform 1 0 144480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1666464484
transform 1 0 152432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1666464484
transform 1 0 160384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1666464484
transform 1 0 168336 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1666464484
transform 1 0 176288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1666464484
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1666464484
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1666464484
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1666464484
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1666464484
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1666464484
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1666464484
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1666464484
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1666464484
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1666464484
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1666464484
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1666464484
transform 1 0 92736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1666464484
transform 1 0 100688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1666464484
transform 1 0 108640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1666464484
transform 1 0 116592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1666464484
transform 1 0 124544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1666464484
transform 1 0 132496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1666464484
transform 1 0 140448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1666464484
transform 1 0 148400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1666464484
transform 1 0 156352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1666464484
transform 1 0 164304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1666464484
transform 1 0 172256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1666464484
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1666464484
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1666464484
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1666464484
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1666464484
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1666464484
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1666464484
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1666464484
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1666464484
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1666464484
transform 1 0 80864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1666464484
transform 1 0 88816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1666464484
transform 1 0 96768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1666464484
transform 1 0 104720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1666464484
transform 1 0 112672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1666464484
transform 1 0 120624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1666464484
transform 1 0 128576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1666464484
transform 1 0 136528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1666464484
transform 1 0 144480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1666464484
transform 1 0 152432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1666464484
transform 1 0 160384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1666464484
transform 1 0 168336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1666464484
transform 1 0 176288 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1666464484
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1666464484
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1666464484
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1666464484
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1666464484
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1666464484
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1666464484
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1666464484
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1666464484
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1666464484
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1666464484
transform 1 0 84784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1666464484
transform 1 0 92736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1666464484
transform 1 0 100688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1666464484
transform 1 0 108640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1666464484
transform 1 0 116592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1666464484
transform 1 0 124544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1666464484
transform 1 0 132496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1666464484
transform 1 0 140448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1666464484
transform 1 0 148400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1666464484
transform 1 0 156352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1666464484
transform 1 0 164304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1666464484
transform 1 0 172256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1666464484
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1666464484
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1666464484
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1666464484
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1666464484
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1666464484
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1666464484
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1666464484
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1666464484
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1666464484
transform 1 0 80864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1666464484
transform 1 0 88816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1666464484
transform 1 0 96768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1666464484
transform 1 0 104720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1666464484
transform 1 0 112672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1666464484
transform 1 0 120624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1666464484
transform 1 0 128576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1666464484
transform 1 0 136528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1666464484
transform 1 0 144480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1666464484
transform 1 0 152432 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1666464484
transform 1 0 160384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1666464484
transform 1 0 168336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1666464484
transform 1 0 176288 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1666464484
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1666464484
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1666464484
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1666464484
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1666464484
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1666464484
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1666464484
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1666464484
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1666464484
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1666464484
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1666464484
transform 1 0 84784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1666464484
transform 1 0 92736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1666464484
transform 1 0 100688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_898
timestamp 1666464484
transform 1 0 108640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_899
timestamp 1666464484
transform 1 0 116592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_900
timestamp 1666464484
transform 1 0 124544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_901
timestamp 1666464484
transform 1 0 132496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_902
timestamp 1666464484
transform 1 0 140448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_903
timestamp 1666464484
transform 1 0 148400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_904
timestamp 1666464484
transform 1 0 156352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_905
timestamp 1666464484
transform 1 0 164304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_906
timestamp 1666464484
transform 1 0 172256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_907
timestamp 1666464484
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_908
timestamp 1666464484
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_909
timestamp 1666464484
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_910
timestamp 1666464484
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_911
timestamp 1666464484
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_912
timestamp 1666464484
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_913
timestamp 1666464484
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_914
timestamp 1666464484
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_915
timestamp 1666464484
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_916
timestamp 1666464484
transform 1 0 80864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_917
timestamp 1666464484
transform 1 0 88816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_918
timestamp 1666464484
transform 1 0 96768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_919
timestamp 1666464484
transform 1 0 104720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_920
timestamp 1666464484
transform 1 0 112672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_921
timestamp 1666464484
transform 1 0 120624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_922
timestamp 1666464484
transform 1 0 128576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_923
timestamp 1666464484
transform 1 0 136528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_924
timestamp 1666464484
transform 1 0 144480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_925
timestamp 1666464484
transform 1 0 152432 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_926
timestamp 1666464484
transform 1 0 160384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_927
timestamp 1666464484
transform 1 0 168336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_928
timestamp 1666464484
transform 1 0 176288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_929
timestamp 1666464484
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_930
timestamp 1666464484
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_931
timestamp 1666464484
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_932
timestamp 1666464484
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_933
timestamp 1666464484
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_934
timestamp 1666464484
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_935
timestamp 1666464484
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_936
timestamp 1666464484
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_937
timestamp 1666464484
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_938
timestamp 1666464484
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_939
timestamp 1666464484
transform 1 0 84784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_940
timestamp 1666464484
transform 1 0 92736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_941
timestamp 1666464484
transform 1 0 100688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_942
timestamp 1666464484
transform 1 0 108640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_943
timestamp 1666464484
transform 1 0 116592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_944
timestamp 1666464484
transform 1 0 124544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_945
timestamp 1666464484
transform 1 0 132496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_946
timestamp 1666464484
transform 1 0 140448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_947
timestamp 1666464484
transform 1 0 148400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_948
timestamp 1666464484
transform 1 0 156352 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_949
timestamp 1666464484
transform 1 0 164304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_950
timestamp 1666464484
transform 1 0 172256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_951
timestamp 1666464484
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_952
timestamp 1666464484
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_953
timestamp 1666464484
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_954
timestamp 1666464484
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_955
timestamp 1666464484
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_956
timestamp 1666464484
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_957
timestamp 1666464484
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_958
timestamp 1666464484
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_959
timestamp 1666464484
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_960
timestamp 1666464484
transform 1 0 80864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_961
timestamp 1666464484
transform 1 0 88816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_962
timestamp 1666464484
transform 1 0 96768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_963
timestamp 1666464484
transform 1 0 104720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_964
timestamp 1666464484
transform 1 0 112672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_965
timestamp 1666464484
transform 1 0 120624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_966
timestamp 1666464484
transform 1 0 128576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_967
timestamp 1666464484
transform 1 0 136528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_968
timestamp 1666464484
transform 1 0 144480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_969
timestamp 1666464484
transform 1 0 152432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_970
timestamp 1666464484
transform 1 0 160384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_971
timestamp 1666464484
transform 1 0 168336 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_972
timestamp 1666464484
transform 1 0 176288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_973
timestamp 1666464484
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_974
timestamp 1666464484
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_975
timestamp 1666464484
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_976
timestamp 1666464484
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_977
timestamp 1666464484
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_978
timestamp 1666464484
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_979
timestamp 1666464484
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_980
timestamp 1666464484
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_981
timestamp 1666464484
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_982
timestamp 1666464484
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_983
timestamp 1666464484
transform 1 0 84784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_984
timestamp 1666464484
transform 1 0 92736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_985
timestamp 1666464484
transform 1 0 100688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_986
timestamp 1666464484
transform 1 0 108640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_987
timestamp 1666464484
transform 1 0 116592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_988
timestamp 1666464484
transform 1 0 124544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_989
timestamp 1666464484
transform 1 0 132496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_990
timestamp 1666464484
transform 1 0 140448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_991
timestamp 1666464484
transform 1 0 148400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_992
timestamp 1666464484
transform 1 0 156352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_993
timestamp 1666464484
transform 1 0 164304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_994
timestamp 1666464484
transform 1 0 172256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_995
timestamp 1666464484
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_996
timestamp 1666464484
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_997
timestamp 1666464484
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_998
timestamp 1666464484
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_999
timestamp 1666464484
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1000
timestamp 1666464484
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1001
timestamp 1666464484
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1002
timestamp 1666464484
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1003
timestamp 1666464484
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1004
timestamp 1666464484
transform 1 0 80864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1005
timestamp 1666464484
transform 1 0 88816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1006
timestamp 1666464484
transform 1 0 96768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1007
timestamp 1666464484
transform 1 0 104720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1008
timestamp 1666464484
transform 1 0 112672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1009
timestamp 1666464484
transform 1 0 120624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1010
timestamp 1666464484
transform 1 0 128576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1011
timestamp 1666464484
transform 1 0 136528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1012
timestamp 1666464484
transform 1 0 144480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1013
timestamp 1666464484
transform 1 0 152432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1014
timestamp 1666464484
transform 1 0 160384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1015
timestamp 1666464484
transform 1 0 168336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1016
timestamp 1666464484
transform 1 0 176288 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1017
timestamp 1666464484
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1018
timestamp 1666464484
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1019
timestamp 1666464484
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1020
timestamp 1666464484
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1021
timestamp 1666464484
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1022
timestamp 1666464484
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1023
timestamp 1666464484
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1024
timestamp 1666464484
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1025
timestamp 1666464484
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1026
timestamp 1666464484
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1027
timestamp 1666464484
transform 1 0 84784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1028
timestamp 1666464484
transform 1 0 92736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1029
timestamp 1666464484
transform 1 0 100688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1030
timestamp 1666464484
transform 1 0 108640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1031
timestamp 1666464484
transform 1 0 116592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1032
timestamp 1666464484
transform 1 0 124544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1033
timestamp 1666464484
transform 1 0 132496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1034
timestamp 1666464484
transform 1 0 140448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1035
timestamp 1666464484
transform 1 0 148400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1036
timestamp 1666464484
transform 1 0 156352 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1037
timestamp 1666464484
transform 1 0 164304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1038
timestamp 1666464484
transform 1 0 172256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1039
timestamp 1666464484
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1040
timestamp 1666464484
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1041
timestamp 1666464484
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1042
timestamp 1666464484
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1043
timestamp 1666464484
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1044
timestamp 1666464484
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1045
timestamp 1666464484
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1046
timestamp 1666464484
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1047
timestamp 1666464484
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1048
timestamp 1666464484
transform 1 0 80864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1049
timestamp 1666464484
transform 1 0 88816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1050
timestamp 1666464484
transform 1 0 96768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1051
timestamp 1666464484
transform 1 0 104720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1052
timestamp 1666464484
transform 1 0 112672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1053
timestamp 1666464484
transform 1 0 120624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1054
timestamp 1666464484
transform 1 0 128576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1055
timestamp 1666464484
transform 1 0 136528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1056
timestamp 1666464484
transform 1 0 144480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1057
timestamp 1666464484
transform 1 0 152432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1058
timestamp 1666464484
transform 1 0 160384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1059
timestamp 1666464484
transform 1 0 168336 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1060
timestamp 1666464484
transform 1 0 176288 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1061
timestamp 1666464484
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1062
timestamp 1666464484
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1063
timestamp 1666464484
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1064
timestamp 1666464484
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1065
timestamp 1666464484
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1066
timestamp 1666464484
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1067
timestamp 1666464484
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1068
timestamp 1666464484
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1069
timestamp 1666464484
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1070
timestamp 1666464484
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1071
timestamp 1666464484
transform 1 0 84784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1072
timestamp 1666464484
transform 1 0 92736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1073
timestamp 1666464484
transform 1 0 100688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1074
timestamp 1666464484
transform 1 0 108640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1075
timestamp 1666464484
transform 1 0 116592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1076
timestamp 1666464484
transform 1 0 124544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1077
timestamp 1666464484
transform 1 0 132496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1078
timestamp 1666464484
transform 1 0 140448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1079
timestamp 1666464484
transform 1 0 148400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1080
timestamp 1666464484
transform 1 0 156352 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1081
timestamp 1666464484
transform 1 0 164304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1082
timestamp 1666464484
transform 1 0 172256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1083
timestamp 1666464484
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1084
timestamp 1666464484
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1085
timestamp 1666464484
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1086
timestamp 1666464484
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1087
timestamp 1666464484
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1088
timestamp 1666464484
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1089
timestamp 1666464484
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1090
timestamp 1666464484
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1091
timestamp 1666464484
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1092
timestamp 1666464484
transform 1 0 80864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1093
timestamp 1666464484
transform 1 0 88816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1094
timestamp 1666464484
transform 1 0 96768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1095
timestamp 1666464484
transform 1 0 104720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1096
timestamp 1666464484
transform 1 0 112672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1097
timestamp 1666464484
transform 1 0 120624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1098
timestamp 1666464484
transform 1 0 128576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1099
timestamp 1666464484
transform 1 0 136528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1100
timestamp 1666464484
transform 1 0 144480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1101
timestamp 1666464484
transform 1 0 152432 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1102
timestamp 1666464484
transform 1 0 160384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1103
timestamp 1666464484
transform 1 0 168336 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1104
timestamp 1666464484
transform 1 0 176288 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1105
timestamp 1666464484
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1106
timestamp 1666464484
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1107
timestamp 1666464484
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1108
timestamp 1666464484
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1109
timestamp 1666464484
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1110
timestamp 1666464484
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1111
timestamp 1666464484
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1112
timestamp 1666464484
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1113
timestamp 1666464484
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1114
timestamp 1666464484
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1115
timestamp 1666464484
transform 1 0 84784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1116
timestamp 1666464484
transform 1 0 92736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1117
timestamp 1666464484
transform 1 0 100688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1118
timestamp 1666464484
transform 1 0 108640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1119
timestamp 1666464484
transform 1 0 116592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1120
timestamp 1666464484
transform 1 0 124544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1121
timestamp 1666464484
transform 1 0 132496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1122
timestamp 1666464484
transform 1 0 140448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1123
timestamp 1666464484
transform 1 0 148400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1124
timestamp 1666464484
transform 1 0 156352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1125
timestamp 1666464484
transform 1 0 164304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1126
timestamp 1666464484
transform 1 0 172256 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1127
timestamp 1666464484
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1128
timestamp 1666464484
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1129
timestamp 1666464484
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1130
timestamp 1666464484
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1131
timestamp 1666464484
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1132
timestamp 1666464484
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1133
timestamp 1666464484
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1134
timestamp 1666464484
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1135
timestamp 1666464484
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1136
timestamp 1666464484
transform 1 0 80864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1137
timestamp 1666464484
transform 1 0 88816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1138
timestamp 1666464484
transform 1 0 96768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1139
timestamp 1666464484
transform 1 0 104720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1140
timestamp 1666464484
transform 1 0 112672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1141
timestamp 1666464484
transform 1 0 120624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1142
timestamp 1666464484
transform 1 0 128576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1143
timestamp 1666464484
transform 1 0 136528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1144
timestamp 1666464484
transform 1 0 144480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1145
timestamp 1666464484
transform 1 0 152432 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1146
timestamp 1666464484
transform 1 0 160384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1147
timestamp 1666464484
transform 1 0 168336 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1148
timestamp 1666464484
transform 1 0 176288 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1149
timestamp 1666464484
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1150
timestamp 1666464484
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1151
timestamp 1666464484
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1152
timestamp 1666464484
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1153
timestamp 1666464484
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1154
timestamp 1666464484
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1155
timestamp 1666464484
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1156
timestamp 1666464484
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1157
timestamp 1666464484
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1158
timestamp 1666464484
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1159
timestamp 1666464484
transform 1 0 84784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1160
timestamp 1666464484
transform 1 0 92736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1161
timestamp 1666464484
transform 1 0 100688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1162
timestamp 1666464484
transform 1 0 108640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1163
timestamp 1666464484
transform 1 0 116592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1164
timestamp 1666464484
transform 1 0 124544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1165
timestamp 1666464484
transform 1 0 132496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1166
timestamp 1666464484
transform 1 0 140448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1167
timestamp 1666464484
transform 1 0 148400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1168
timestamp 1666464484
transform 1 0 156352 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1169
timestamp 1666464484
transform 1 0 164304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1170
timestamp 1666464484
transform 1 0 172256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1171
timestamp 1666464484
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1172
timestamp 1666464484
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1173
timestamp 1666464484
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1174
timestamp 1666464484
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1175
timestamp 1666464484
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1176
timestamp 1666464484
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1177
timestamp 1666464484
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1178
timestamp 1666464484
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1179
timestamp 1666464484
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1180
timestamp 1666464484
transform 1 0 80864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1181
timestamp 1666464484
transform 1 0 88816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1182
timestamp 1666464484
transform 1 0 96768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1183
timestamp 1666464484
transform 1 0 104720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1184
timestamp 1666464484
transform 1 0 112672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1185
timestamp 1666464484
transform 1 0 120624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1186
timestamp 1666464484
transform 1 0 128576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1187
timestamp 1666464484
transform 1 0 136528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1188
timestamp 1666464484
transform 1 0 144480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1189
timestamp 1666464484
transform 1 0 152432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1190
timestamp 1666464484
transform 1 0 160384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1191
timestamp 1666464484
transform 1 0 168336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1192
timestamp 1666464484
transform 1 0 176288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1193
timestamp 1666464484
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1194
timestamp 1666464484
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1195
timestamp 1666464484
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1196
timestamp 1666464484
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1197
timestamp 1666464484
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1198
timestamp 1666464484
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1199
timestamp 1666464484
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1200
timestamp 1666464484
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1201
timestamp 1666464484
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1202
timestamp 1666464484
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1203
timestamp 1666464484
transform 1 0 84784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1204
timestamp 1666464484
transform 1 0 92736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1205
timestamp 1666464484
transform 1 0 100688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1206
timestamp 1666464484
transform 1 0 108640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1207
timestamp 1666464484
transform 1 0 116592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1208
timestamp 1666464484
transform 1 0 124544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1209
timestamp 1666464484
transform 1 0 132496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1210
timestamp 1666464484
transform 1 0 140448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1211
timestamp 1666464484
transform 1 0 148400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1212
timestamp 1666464484
transform 1 0 156352 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1213
timestamp 1666464484
transform 1 0 164304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1214
timestamp 1666464484
transform 1 0 172256 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1215
timestamp 1666464484
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1216
timestamp 1666464484
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1217
timestamp 1666464484
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1218
timestamp 1666464484
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1219
timestamp 1666464484
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1220
timestamp 1666464484
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1221
timestamp 1666464484
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1222
timestamp 1666464484
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1223
timestamp 1666464484
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1224
timestamp 1666464484
transform 1 0 80864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1225
timestamp 1666464484
transform 1 0 88816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1226
timestamp 1666464484
transform 1 0 96768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1227
timestamp 1666464484
transform 1 0 104720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1228
timestamp 1666464484
transform 1 0 112672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1229
timestamp 1666464484
transform 1 0 120624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1230
timestamp 1666464484
transform 1 0 128576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1231
timestamp 1666464484
transform 1 0 136528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1232
timestamp 1666464484
transform 1 0 144480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1233
timestamp 1666464484
transform 1 0 152432 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1234
timestamp 1666464484
transform 1 0 160384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1235
timestamp 1666464484
transform 1 0 168336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1236
timestamp 1666464484
transform 1 0 176288 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1237
timestamp 1666464484
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1238
timestamp 1666464484
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1239
timestamp 1666464484
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1240
timestamp 1666464484
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1241
timestamp 1666464484
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1242
timestamp 1666464484
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1243
timestamp 1666464484
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1244
timestamp 1666464484
transform 1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1245
timestamp 1666464484
transform 1 0 68880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1246
timestamp 1666464484
transform 1 0 76832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1247
timestamp 1666464484
transform 1 0 84784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1248
timestamp 1666464484
transform 1 0 92736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1249
timestamp 1666464484
transform 1 0 100688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1250
timestamp 1666464484
transform 1 0 108640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1251
timestamp 1666464484
transform 1 0 116592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1252
timestamp 1666464484
transform 1 0 124544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1253
timestamp 1666464484
transform 1 0 132496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1254
timestamp 1666464484
transform 1 0 140448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1255
timestamp 1666464484
transform 1 0 148400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1256
timestamp 1666464484
transform 1 0 156352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1257
timestamp 1666464484
transform 1 0 164304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1258
timestamp 1666464484
transform 1 0 172256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1259
timestamp 1666464484
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1260
timestamp 1666464484
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1261
timestamp 1666464484
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1262
timestamp 1666464484
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1263
timestamp 1666464484
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1264
timestamp 1666464484
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1265
timestamp 1666464484
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1266
timestamp 1666464484
transform 1 0 64960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1267
timestamp 1666464484
transform 1 0 72912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1268
timestamp 1666464484
transform 1 0 80864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1269
timestamp 1666464484
transform 1 0 88816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1270
timestamp 1666464484
transform 1 0 96768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1271
timestamp 1666464484
transform 1 0 104720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1272
timestamp 1666464484
transform 1 0 112672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1273
timestamp 1666464484
transform 1 0 120624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1274
timestamp 1666464484
transform 1 0 128576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1275
timestamp 1666464484
transform 1 0 136528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1276
timestamp 1666464484
transform 1 0 144480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1277
timestamp 1666464484
transform 1 0 152432 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1278
timestamp 1666464484
transform 1 0 160384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1279
timestamp 1666464484
transform 1 0 168336 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1280
timestamp 1666464484
transform 1 0 176288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1281
timestamp 1666464484
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1282
timestamp 1666464484
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1283
timestamp 1666464484
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1284
timestamp 1666464484
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1285
timestamp 1666464484
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1286
timestamp 1666464484
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1287
timestamp 1666464484
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1288
timestamp 1666464484
transform 1 0 60928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1289
timestamp 1666464484
transform 1 0 68880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1290
timestamp 1666464484
transform 1 0 76832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1291
timestamp 1666464484
transform 1 0 84784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1292
timestamp 1666464484
transform 1 0 92736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1293
timestamp 1666464484
transform 1 0 100688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1294
timestamp 1666464484
transform 1 0 108640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1295
timestamp 1666464484
transform 1 0 116592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1296
timestamp 1666464484
transform 1 0 124544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1297
timestamp 1666464484
transform 1 0 132496 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1298
timestamp 1666464484
transform 1 0 140448 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1299
timestamp 1666464484
transform 1 0 148400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1300
timestamp 1666464484
transform 1 0 156352 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1301
timestamp 1666464484
transform 1 0 164304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1302
timestamp 1666464484
transform 1 0 172256 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1303
timestamp 1666464484
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1304
timestamp 1666464484
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1305
timestamp 1666464484
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1306
timestamp 1666464484
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1307
timestamp 1666464484
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1308
timestamp 1666464484
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1309
timestamp 1666464484
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1310
timestamp 1666464484
transform 1 0 64960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1311
timestamp 1666464484
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1312
timestamp 1666464484
transform 1 0 80864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1313
timestamp 1666464484
transform 1 0 88816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1314
timestamp 1666464484
transform 1 0 96768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1315
timestamp 1666464484
transform 1 0 104720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1316
timestamp 1666464484
transform 1 0 112672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1317
timestamp 1666464484
transform 1 0 120624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1318
timestamp 1666464484
transform 1 0 128576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1319
timestamp 1666464484
transform 1 0 136528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1320
timestamp 1666464484
transform 1 0 144480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1321
timestamp 1666464484
transform 1 0 152432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1322
timestamp 1666464484
transform 1 0 160384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1323
timestamp 1666464484
transform 1 0 168336 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1324
timestamp 1666464484
transform 1 0 176288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1325
timestamp 1666464484
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1326
timestamp 1666464484
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1327
timestamp 1666464484
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1328
timestamp 1666464484
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1329
timestamp 1666464484
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1330
timestamp 1666464484
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1331
timestamp 1666464484
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1332
timestamp 1666464484
transform 1 0 60928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1333
timestamp 1666464484
transform 1 0 68880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1334
timestamp 1666464484
transform 1 0 76832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1335
timestamp 1666464484
transform 1 0 84784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1336
timestamp 1666464484
transform 1 0 92736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1337
timestamp 1666464484
transform 1 0 100688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1338
timestamp 1666464484
transform 1 0 108640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1339
timestamp 1666464484
transform 1 0 116592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1340
timestamp 1666464484
transform 1 0 124544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1341
timestamp 1666464484
transform 1 0 132496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1342
timestamp 1666464484
transform 1 0 140448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1343
timestamp 1666464484
transform 1 0 148400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1344
timestamp 1666464484
transform 1 0 156352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1345
timestamp 1666464484
transform 1 0 164304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1346
timestamp 1666464484
transform 1 0 172256 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1347
timestamp 1666464484
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1348
timestamp 1666464484
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1349
timestamp 1666464484
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1350
timestamp 1666464484
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1351
timestamp 1666464484
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1352
timestamp 1666464484
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1353
timestamp 1666464484
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1354
timestamp 1666464484
transform 1 0 64960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1355
timestamp 1666464484
transform 1 0 72912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1356
timestamp 1666464484
transform 1 0 80864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1357
timestamp 1666464484
transform 1 0 88816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1358
timestamp 1666464484
transform 1 0 96768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1359
timestamp 1666464484
transform 1 0 104720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1360
timestamp 1666464484
transform 1 0 112672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1361
timestamp 1666464484
transform 1 0 120624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1362
timestamp 1666464484
transform 1 0 128576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1363
timestamp 1666464484
transform 1 0 136528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1364
timestamp 1666464484
transform 1 0 144480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1365
timestamp 1666464484
transform 1 0 152432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1366
timestamp 1666464484
transform 1 0 160384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1367
timestamp 1666464484
transform 1 0 168336 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1368
timestamp 1666464484
transform 1 0 176288 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1369
timestamp 1666464484
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1370
timestamp 1666464484
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1371
timestamp 1666464484
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1372
timestamp 1666464484
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1373
timestamp 1666464484
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1374
timestamp 1666464484
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1375
timestamp 1666464484
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1376
timestamp 1666464484
transform 1 0 60928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1377
timestamp 1666464484
transform 1 0 68880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1378
timestamp 1666464484
transform 1 0 76832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1379
timestamp 1666464484
transform 1 0 84784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1380
timestamp 1666464484
transform 1 0 92736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1381
timestamp 1666464484
transform 1 0 100688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1382
timestamp 1666464484
transform 1 0 108640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1383
timestamp 1666464484
transform 1 0 116592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1384
timestamp 1666464484
transform 1 0 124544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1385
timestamp 1666464484
transform 1 0 132496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1386
timestamp 1666464484
transform 1 0 140448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1387
timestamp 1666464484
transform 1 0 148400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1388
timestamp 1666464484
transform 1 0 156352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1389
timestamp 1666464484
transform 1 0 164304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1390
timestamp 1666464484
transform 1 0 172256 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1391
timestamp 1666464484
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1392
timestamp 1666464484
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1393
timestamp 1666464484
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1394
timestamp 1666464484
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1395
timestamp 1666464484
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1396
timestamp 1666464484
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1397
timestamp 1666464484
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1398
timestamp 1666464484
transform 1 0 64960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1399
timestamp 1666464484
transform 1 0 72912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1400
timestamp 1666464484
transform 1 0 80864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1401
timestamp 1666464484
transform 1 0 88816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1402
timestamp 1666464484
transform 1 0 96768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1403
timestamp 1666464484
transform 1 0 104720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1404
timestamp 1666464484
transform 1 0 112672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1405
timestamp 1666464484
transform 1 0 120624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1406
timestamp 1666464484
transform 1 0 128576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1407
timestamp 1666464484
transform 1 0 136528 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1408
timestamp 1666464484
transform 1 0 144480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1409
timestamp 1666464484
transform 1 0 152432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1410
timestamp 1666464484
transform 1 0 160384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1411
timestamp 1666464484
transform 1 0 168336 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1412
timestamp 1666464484
transform 1 0 176288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1413
timestamp 1666464484
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1414
timestamp 1666464484
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1415
timestamp 1666464484
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1416
timestamp 1666464484
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1417
timestamp 1666464484
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1418
timestamp 1666464484
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1419
timestamp 1666464484
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1420
timestamp 1666464484
transform 1 0 60928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1421
timestamp 1666464484
transform 1 0 68880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1422
timestamp 1666464484
transform 1 0 76832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1423
timestamp 1666464484
transform 1 0 84784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1424
timestamp 1666464484
transform 1 0 92736 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1425
timestamp 1666464484
transform 1 0 100688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1426
timestamp 1666464484
transform 1 0 108640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1427
timestamp 1666464484
transform 1 0 116592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1428
timestamp 1666464484
transform 1 0 124544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1429
timestamp 1666464484
transform 1 0 132496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1430
timestamp 1666464484
transform 1 0 140448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1431
timestamp 1666464484
transform 1 0 148400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1432
timestamp 1666464484
transform 1 0 156352 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1433
timestamp 1666464484
transform 1 0 164304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1434
timestamp 1666464484
transform 1 0 172256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1435
timestamp 1666464484
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1436
timestamp 1666464484
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1437
timestamp 1666464484
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1438
timestamp 1666464484
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1439
timestamp 1666464484
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1440
timestamp 1666464484
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1441
timestamp 1666464484
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1442
timestamp 1666464484
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1443
timestamp 1666464484
transform 1 0 72912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1444
timestamp 1666464484
transform 1 0 80864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1445
timestamp 1666464484
transform 1 0 88816 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1446
timestamp 1666464484
transform 1 0 96768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1447
timestamp 1666464484
transform 1 0 104720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1448
timestamp 1666464484
transform 1 0 112672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1449
timestamp 1666464484
transform 1 0 120624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1450
timestamp 1666464484
transform 1 0 128576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1451
timestamp 1666464484
transform 1 0 136528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1452
timestamp 1666464484
transform 1 0 144480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1453
timestamp 1666464484
transform 1 0 152432 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1454
timestamp 1666464484
transform 1 0 160384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1455
timestamp 1666464484
transform 1 0 168336 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1456
timestamp 1666464484
transform 1 0 176288 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1457
timestamp 1666464484
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1458
timestamp 1666464484
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1459
timestamp 1666464484
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1460
timestamp 1666464484
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1461
timestamp 1666464484
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1462
timestamp 1666464484
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1463
timestamp 1666464484
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1464
timestamp 1666464484
transform 1 0 60928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1465
timestamp 1666464484
transform 1 0 68880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1466
timestamp 1666464484
transform 1 0 76832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1467
timestamp 1666464484
transform 1 0 84784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1468
timestamp 1666464484
transform 1 0 92736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1469
timestamp 1666464484
transform 1 0 100688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1470
timestamp 1666464484
transform 1 0 108640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1471
timestamp 1666464484
transform 1 0 116592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1472
timestamp 1666464484
transform 1 0 124544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1473
timestamp 1666464484
transform 1 0 132496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1474
timestamp 1666464484
transform 1 0 140448 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1475
timestamp 1666464484
transform 1 0 148400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1476
timestamp 1666464484
transform 1 0 156352 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1477
timestamp 1666464484
transform 1 0 164304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1478
timestamp 1666464484
transform 1 0 172256 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1479
timestamp 1666464484
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1480
timestamp 1666464484
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1481
timestamp 1666464484
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1482
timestamp 1666464484
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1483
timestamp 1666464484
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1484
timestamp 1666464484
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1485
timestamp 1666464484
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1486
timestamp 1666464484
transform 1 0 64960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1487
timestamp 1666464484
transform 1 0 72912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1488
timestamp 1666464484
transform 1 0 80864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1489
timestamp 1666464484
transform 1 0 88816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1490
timestamp 1666464484
transform 1 0 96768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1491
timestamp 1666464484
transform 1 0 104720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1492
timestamp 1666464484
transform 1 0 112672 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1493
timestamp 1666464484
transform 1 0 120624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1494
timestamp 1666464484
transform 1 0 128576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1495
timestamp 1666464484
transform 1 0 136528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1496
timestamp 1666464484
transform 1 0 144480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1497
timestamp 1666464484
transform 1 0 152432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1498
timestamp 1666464484
transform 1 0 160384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1499
timestamp 1666464484
transform 1 0 168336 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1500
timestamp 1666464484
transform 1 0 176288 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1501
timestamp 1666464484
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1502
timestamp 1666464484
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1503
timestamp 1666464484
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1504
timestamp 1666464484
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1505
timestamp 1666464484
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1506
timestamp 1666464484
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1507
timestamp 1666464484
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1508
timestamp 1666464484
transform 1 0 60928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1509
timestamp 1666464484
transform 1 0 68880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1510
timestamp 1666464484
transform 1 0 76832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1511
timestamp 1666464484
transform 1 0 84784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1512
timestamp 1666464484
transform 1 0 92736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1513
timestamp 1666464484
transform 1 0 100688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1514
timestamp 1666464484
transform 1 0 108640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1515
timestamp 1666464484
transform 1 0 116592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1516
timestamp 1666464484
transform 1 0 124544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1517
timestamp 1666464484
transform 1 0 132496 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1518
timestamp 1666464484
transform 1 0 140448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1519
timestamp 1666464484
transform 1 0 148400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1520
timestamp 1666464484
transform 1 0 156352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1521
timestamp 1666464484
transform 1 0 164304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1522
timestamp 1666464484
transform 1 0 172256 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1523
timestamp 1666464484
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1524
timestamp 1666464484
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1525
timestamp 1666464484
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1526
timestamp 1666464484
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1527
timestamp 1666464484
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1528
timestamp 1666464484
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1529
timestamp 1666464484
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1530
timestamp 1666464484
transform 1 0 64960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1531
timestamp 1666464484
transform 1 0 72912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1532
timestamp 1666464484
transform 1 0 80864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1533
timestamp 1666464484
transform 1 0 88816 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1534
timestamp 1666464484
transform 1 0 96768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1535
timestamp 1666464484
transform 1 0 104720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1536
timestamp 1666464484
transform 1 0 112672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1537
timestamp 1666464484
transform 1 0 120624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1538
timestamp 1666464484
transform 1 0 128576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1539
timestamp 1666464484
transform 1 0 136528 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1540
timestamp 1666464484
transform 1 0 144480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1541
timestamp 1666464484
transform 1 0 152432 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1542
timestamp 1666464484
transform 1 0 160384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1543
timestamp 1666464484
transform 1 0 168336 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1544
timestamp 1666464484
transform 1 0 176288 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1545
timestamp 1666464484
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1546
timestamp 1666464484
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1547
timestamp 1666464484
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1548
timestamp 1666464484
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1549
timestamp 1666464484
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1550
timestamp 1666464484
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1551
timestamp 1666464484
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1552
timestamp 1666464484
transform 1 0 60928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1553
timestamp 1666464484
transform 1 0 68880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1554
timestamp 1666464484
transform 1 0 76832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1555
timestamp 1666464484
transform 1 0 84784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1556
timestamp 1666464484
transform 1 0 92736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1557
timestamp 1666464484
transform 1 0 100688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1558
timestamp 1666464484
transform 1 0 108640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1559
timestamp 1666464484
transform 1 0 116592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1560
timestamp 1666464484
transform 1 0 124544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1561
timestamp 1666464484
transform 1 0 132496 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1562
timestamp 1666464484
transform 1 0 140448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1563
timestamp 1666464484
transform 1 0 148400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1564
timestamp 1666464484
transform 1 0 156352 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1565
timestamp 1666464484
transform 1 0 164304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1566
timestamp 1666464484
transform 1 0 172256 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1567
timestamp 1666464484
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1568
timestamp 1666464484
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1569
timestamp 1666464484
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1570
timestamp 1666464484
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1571
timestamp 1666464484
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1572
timestamp 1666464484
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1573
timestamp 1666464484
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1574
timestamp 1666464484
transform 1 0 64960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1575
timestamp 1666464484
transform 1 0 72912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1576
timestamp 1666464484
transform 1 0 80864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1577
timestamp 1666464484
transform 1 0 88816 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1578
timestamp 1666464484
transform 1 0 96768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1579
timestamp 1666464484
transform 1 0 104720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1580
timestamp 1666464484
transform 1 0 112672 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1581
timestamp 1666464484
transform 1 0 120624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1582
timestamp 1666464484
transform 1 0 128576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1583
timestamp 1666464484
transform 1 0 136528 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1584
timestamp 1666464484
transform 1 0 144480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1585
timestamp 1666464484
transform 1 0 152432 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1586
timestamp 1666464484
transform 1 0 160384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1587
timestamp 1666464484
transform 1 0 168336 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1588
timestamp 1666464484
transform 1 0 176288 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1589
timestamp 1666464484
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1590
timestamp 1666464484
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1591
timestamp 1666464484
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1592
timestamp 1666464484
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1593
timestamp 1666464484
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1594
timestamp 1666464484
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1595
timestamp 1666464484
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1596
timestamp 1666464484
transform 1 0 60928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1597
timestamp 1666464484
transform 1 0 68880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1598
timestamp 1666464484
transform 1 0 76832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1599
timestamp 1666464484
transform 1 0 84784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1600
timestamp 1666464484
transform 1 0 92736 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1601
timestamp 1666464484
transform 1 0 100688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1602
timestamp 1666464484
transform 1 0 108640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1603
timestamp 1666464484
transform 1 0 116592 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1604
timestamp 1666464484
transform 1 0 124544 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1605
timestamp 1666464484
transform 1 0 132496 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1606
timestamp 1666464484
transform 1 0 140448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1607
timestamp 1666464484
transform 1 0 148400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1608
timestamp 1666464484
transform 1 0 156352 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1609
timestamp 1666464484
transform 1 0 164304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1610
timestamp 1666464484
transform 1 0 172256 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1611
timestamp 1666464484
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1612
timestamp 1666464484
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1613
timestamp 1666464484
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1614
timestamp 1666464484
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1615
timestamp 1666464484
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1616
timestamp 1666464484
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1617
timestamp 1666464484
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1618
timestamp 1666464484
transform 1 0 64960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1619
timestamp 1666464484
transform 1 0 72912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1620
timestamp 1666464484
transform 1 0 80864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1621
timestamp 1666464484
transform 1 0 88816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1622
timestamp 1666464484
transform 1 0 96768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1623
timestamp 1666464484
transform 1 0 104720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1624
timestamp 1666464484
transform 1 0 112672 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1625
timestamp 1666464484
transform 1 0 120624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1626
timestamp 1666464484
transform 1 0 128576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1627
timestamp 1666464484
transform 1 0 136528 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1628
timestamp 1666464484
transform 1 0 144480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1629
timestamp 1666464484
transform 1 0 152432 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1630
timestamp 1666464484
transform 1 0 160384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1631
timestamp 1666464484
transform 1 0 168336 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1632
timestamp 1666464484
transform 1 0 176288 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1633
timestamp 1666464484
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1634
timestamp 1666464484
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1635
timestamp 1666464484
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1636
timestamp 1666464484
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1637
timestamp 1666464484
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1638
timestamp 1666464484
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1639
timestamp 1666464484
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1640
timestamp 1666464484
transform 1 0 60928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1641
timestamp 1666464484
transform 1 0 68880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1642
timestamp 1666464484
transform 1 0 76832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1643
timestamp 1666464484
transform 1 0 84784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1644
timestamp 1666464484
transform 1 0 92736 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1645
timestamp 1666464484
transform 1 0 100688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1646
timestamp 1666464484
transform 1 0 108640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1647
timestamp 1666464484
transform 1 0 116592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1648
timestamp 1666464484
transform 1 0 124544 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1649
timestamp 1666464484
transform 1 0 132496 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1650
timestamp 1666464484
transform 1 0 140448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1651
timestamp 1666464484
transform 1 0 148400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1652
timestamp 1666464484
transform 1 0 156352 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1653
timestamp 1666464484
transform 1 0 164304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1654
timestamp 1666464484
transform 1 0 172256 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1655
timestamp 1666464484
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1656
timestamp 1666464484
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1657
timestamp 1666464484
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1658
timestamp 1666464484
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1659
timestamp 1666464484
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1660
timestamp 1666464484
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1661
timestamp 1666464484
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1662
timestamp 1666464484
transform 1 0 64960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1663
timestamp 1666464484
transform 1 0 72912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1664
timestamp 1666464484
transform 1 0 80864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1665
timestamp 1666464484
transform 1 0 88816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1666
timestamp 1666464484
transform 1 0 96768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1667
timestamp 1666464484
transform 1 0 104720 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1668
timestamp 1666464484
transform 1 0 112672 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1669
timestamp 1666464484
transform 1 0 120624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1670
timestamp 1666464484
transform 1 0 128576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1671
timestamp 1666464484
transform 1 0 136528 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1672
timestamp 1666464484
transform 1 0 144480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1673
timestamp 1666464484
transform 1 0 152432 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1674
timestamp 1666464484
transform 1 0 160384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1675
timestamp 1666464484
transform 1 0 168336 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1676
timestamp 1666464484
transform 1 0 176288 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1677
timestamp 1666464484
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1678
timestamp 1666464484
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1679
timestamp 1666464484
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1680
timestamp 1666464484
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1681
timestamp 1666464484
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1682
timestamp 1666464484
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1683
timestamp 1666464484
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1684
timestamp 1666464484
transform 1 0 60928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1685
timestamp 1666464484
transform 1 0 68880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1686
timestamp 1666464484
transform 1 0 76832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1687
timestamp 1666464484
transform 1 0 84784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1688
timestamp 1666464484
transform 1 0 92736 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1689
timestamp 1666464484
transform 1 0 100688 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1690
timestamp 1666464484
transform 1 0 108640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1691
timestamp 1666464484
transform 1 0 116592 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1692
timestamp 1666464484
transform 1 0 124544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1693
timestamp 1666464484
transform 1 0 132496 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1694
timestamp 1666464484
transform 1 0 140448 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1695
timestamp 1666464484
transform 1 0 148400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1696
timestamp 1666464484
transform 1 0 156352 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1697
timestamp 1666464484
transform 1 0 164304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1698
timestamp 1666464484
transform 1 0 172256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1699
timestamp 1666464484
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1700
timestamp 1666464484
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1701
timestamp 1666464484
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1702
timestamp 1666464484
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1703
timestamp 1666464484
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1704
timestamp 1666464484
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1705
timestamp 1666464484
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1706
timestamp 1666464484
transform 1 0 64960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1707
timestamp 1666464484
transform 1 0 72912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1708
timestamp 1666464484
transform 1 0 80864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1709
timestamp 1666464484
transform 1 0 88816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1710
timestamp 1666464484
transform 1 0 96768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1711
timestamp 1666464484
transform 1 0 104720 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1712
timestamp 1666464484
transform 1 0 112672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1713
timestamp 1666464484
transform 1 0 120624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1714
timestamp 1666464484
transform 1 0 128576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1715
timestamp 1666464484
transform 1 0 136528 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1716
timestamp 1666464484
transform 1 0 144480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1717
timestamp 1666464484
transform 1 0 152432 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1718
timestamp 1666464484
transform 1 0 160384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1719
timestamp 1666464484
transform 1 0 168336 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1720
timestamp 1666464484
transform 1 0 176288 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1721
timestamp 1666464484
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1722
timestamp 1666464484
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1723
timestamp 1666464484
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1724
timestamp 1666464484
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1725
timestamp 1666464484
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1726
timestamp 1666464484
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1727
timestamp 1666464484
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1728
timestamp 1666464484
transform 1 0 60928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1729
timestamp 1666464484
transform 1 0 68880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1730
timestamp 1666464484
transform 1 0 76832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1731
timestamp 1666464484
transform 1 0 84784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1732
timestamp 1666464484
transform 1 0 92736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1733
timestamp 1666464484
transform 1 0 100688 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1734
timestamp 1666464484
transform 1 0 108640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1735
timestamp 1666464484
transform 1 0 116592 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1736
timestamp 1666464484
transform 1 0 124544 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1737
timestamp 1666464484
transform 1 0 132496 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1738
timestamp 1666464484
transform 1 0 140448 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1739
timestamp 1666464484
transform 1 0 148400 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1740
timestamp 1666464484
transform 1 0 156352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1741
timestamp 1666464484
transform 1 0 164304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1742
timestamp 1666464484
transform 1 0 172256 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1743
timestamp 1666464484
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1744
timestamp 1666464484
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1745
timestamp 1666464484
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1746
timestamp 1666464484
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1747
timestamp 1666464484
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1748
timestamp 1666464484
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1749
timestamp 1666464484
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1750
timestamp 1666464484
transform 1 0 64960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1751
timestamp 1666464484
transform 1 0 72912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1752
timestamp 1666464484
transform 1 0 80864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1753
timestamp 1666464484
transform 1 0 88816 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1754
timestamp 1666464484
transform 1 0 96768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1755
timestamp 1666464484
transform 1 0 104720 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1756
timestamp 1666464484
transform 1 0 112672 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1757
timestamp 1666464484
transform 1 0 120624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1758
timestamp 1666464484
transform 1 0 128576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1759
timestamp 1666464484
transform 1 0 136528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1760
timestamp 1666464484
transform 1 0 144480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1761
timestamp 1666464484
transform 1 0 152432 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1762
timestamp 1666464484
transform 1 0 160384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1763
timestamp 1666464484
transform 1 0 168336 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1764
timestamp 1666464484
transform 1 0 176288 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1765
timestamp 1666464484
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1766
timestamp 1666464484
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1767
timestamp 1666464484
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1768
timestamp 1666464484
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1769
timestamp 1666464484
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1770
timestamp 1666464484
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1771
timestamp 1666464484
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1772
timestamp 1666464484
transform 1 0 60928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1773
timestamp 1666464484
transform 1 0 68880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1774
timestamp 1666464484
transform 1 0 76832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1775
timestamp 1666464484
transform 1 0 84784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1776
timestamp 1666464484
transform 1 0 92736 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1777
timestamp 1666464484
transform 1 0 100688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1778
timestamp 1666464484
transform 1 0 108640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1779
timestamp 1666464484
transform 1 0 116592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1780
timestamp 1666464484
transform 1 0 124544 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1781
timestamp 1666464484
transform 1 0 132496 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1782
timestamp 1666464484
transform 1 0 140448 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1783
timestamp 1666464484
transform 1 0 148400 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1784
timestamp 1666464484
transform 1 0 156352 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1785
timestamp 1666464484
transform 1 0 164304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1786
timestamp 1666464484
transform 1 0 172256 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1787
timestamp 1666464484
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1788
timestamp 1666464484
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1789
timestamp 1666464484
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1790
timestamp 1666464484
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1791
timestamp 1666464484
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1792
timestamp 1666464484
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1793
timestamp 1666464484
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1794
timestamp 1666464484
transform 1 0 64960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1795
timestamp 1666464484
transform 1 0 72912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1796
timestamp 1666464484
transform 1 0 80864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1797
timestamp 1666464484
transform 1 0 88816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1798
timestamp 1666464484
transform 1 0 96768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1799
timestamp 1666464484
transform 1 0 104720 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1800
timestamp 1666464484
transform 1 0 112672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1801
timestamp 1666464484
transform 1 0 120624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1802
timestamp 1666464484
transform 1 0 128576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1803
timestamp 1666464484
transform 1 0 136528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1804
timestamp 1666464484
transform 1 0 144480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1805
timestamp 1666464484
transform 1 0 152432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1806
timestamp 1666464484
transform 1 0 160384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1807
timestamp 1666464484
transform 1 0 168336 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1808
timestamp 1666464484
transform 1 0 176288 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1809
timestamp 1666464484
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1810
timestamp 1666464484
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1811
timestamp 1666464484
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1812
timestamp 1666464484
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1813
timestamp 1666464484
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1814
timestamp 1666464484
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1815
timestamp 1666464484
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1816
timestamp 1666464484
transform 1 0 60928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1817
timestamp 1666464484
transform 1 0 68880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1818
timestamp 1666464484
transform 1 0 76832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1819
timestamp 1666464484
transform 1 0 84784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1820
timestamp 1666464484
transform 1 0 92736 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1821
timestamp 1666464484
transform 1 0 100688 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1822
timestamp 1666464484
transform 1 0 108640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1823
timestamp 1666464484
transform 1 0 116592 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1824
timestamp 1666464484
transform 1 0 124544 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1825
timestamp 1666464484
transform 1 0 132496 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1826
timestamp 1666464484
transform 1 0 140448 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1827
timestamp 1666464484
transform 1 0 148400 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1828
timestamp 1666464484
transform 1 0 156352 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1829
timestamp 1666464484
transform 1 0 164304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1830
timestamp 1666464484
transform 1 0 172256 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1831
timestamp 1666464484
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1832
timestamp 1666464484
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1833
timestamp 1666464484
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1834
timestamp 1666464484
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1835
timestamp 1666464484
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1836
timestamp 1666464484
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1837
timestamp 1666464484
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1838
timestamp 1666464484
transform 1 0 64960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1839
timestamp 1666464484
transform 1 0 72912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1840
timestamp 1666464484
transform 1 0 80864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1841
timestamp 1666464484
transform 1 0 88816 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1842
timestamp 1666464484
transform 1 0 96768 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1843
timestamp 1666464484
transform 1 0 104720 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1844
timestamp 1666464484
transform 1 0 112672 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1845
timestamp 1666464484
transform 1 0 120624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1846
timestamp 1666464484
transform 1 0 128576 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1847
timestamp 1666464484
transform 1 0 136528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1848
timestamp 1666464484
transform 1 0 144480 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1849
timestamp 1666464484
transform 1 0 152432 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1850
timestamp 1666464484
transform 1 0 160384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1851
timestamp 1666464484
transform 1 0 168336 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1852
timestamp 1666464484
transform 1 0 176288 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1853
timestamp 1666464484
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1854
timestamp 1666464484
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1855
timestamp 1666464484
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1856
timestamp 1666464484
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1857
timestamp 1666464484
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1858
timestamp 1666464484
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1859
timestamp 1666464484
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1860
timestamp 1666464484
transform 1 0 60928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1861
timestamp 1666464484
transform 1 0 68880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1862
timestamp 1666464484
transform 1 0 76832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1863
timestamp 1666464484
transform 1 0 84784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1864
timestamp 1666464484
transform 1 0 92736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1865
timestamp 1666464484
transform 1 0 100688 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1866
timestamp 1666464484
transform 1 0 108640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1867
timestamp 1666464484
transform 1 0 116592 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1868
timestamp 1666464484
transform 1 0 124544 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1869
timestamp 1666464484
transform 1 0 132496 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1870
timestamp 1666464484
transform 1 0 140448 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1871
timestamp 1666464484
transform 1 0 148400 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1872
timestamp 1666464484
transform 1 0 156352 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1873
timestamp 1666464484
transform 1 0 164304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1874
timestamp 1666464484
transform 1 0 172256 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1875
timestamp 1666464484
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1876
timestamp 1666464484
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1877
timestamp 1666464484
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1878
timestamp 1666464484
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1879
timestamp 1666464484
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1880
timestamp 1666464484
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1881
timestamp 1666464484
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1882
timestamp 1666464484
transform 1 0 64960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1883
timestamp 1666464484
transform 1 0 72912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1884
timestamp 1666464484
transform 1 0 80864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1885
timestamp 1666464484
transform 1 0 88816 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1886
timestamp 1666464484
transform 1 0 96768 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1887
timestamp 1666464484
transform 1 0 104720 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1888
timestamp 1666464484
transform 1 0 112672 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1889
timestamp 1666464484
transform 1 0 120624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1890
timestamp 1666464484
transform 1 0 128576 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1891
timestamp 1666464484
transform 1 0 136528 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1892
timestamp 1666464484
transform 1 0 144480 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1893
timestamp 1666464484
transform 1 0 152432 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1894
timestamp 1666464484
transform 1 0 160384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1895
timestamp 1666464484
transform 1 0 168336 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1896
timestamp 1666464484
transform 1 0 176288 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1897
timestamp 1666464484
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1898
timestamp 1666464484
transform 1 0 13216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1899
timestamp 1666464484
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1900
timestamp 1666464484
transform 1 0 29120 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1901
timestamp 1666464484
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1902
timestamp 1666464484
transform 1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1903
timestamp 1666464484
transform 1 0 52976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1904
timestamp 1666464484
transform 1 0 60928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1905
timestamp 1666464484
transform 1 0 68880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1906
timestamp 1666464484
transform 1 0 76832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1907
timestamp 1666464484
transform 1 0 84784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1908
timestamp 1666464484
transform 1 0 92736 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1909
timestamp 1666464484
transform 1 0 100688 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1910
timestamp 1666464484
transform 1 0 108640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1911
timestamp 1666464484
transform 1 0 116592 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1912
timestamp 1666464484
transform 1 0 124544 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1913
timestamp 1666464484
transform 1 0 132496 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1914
timestamp 1666464484
transform 1 0 140448 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1915
timestamp 1666464484
transform 1 0 148400 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1916
timestamp 1666464484
transform 1 0 156352 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1917
timestamp 1666464484
transform 1 0 164304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1918
timestamp 1666464484
transform 1 0 172256 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1919
timestamp 1666464484
transform 1 0 9296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1920
timestamp 1666464484
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1921
timestamp 1666464484
transform 1 0 25200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1922
timestamp 1666464484
transform 1 0 33152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1923
timestamp 1666464484
transform 1 0 41104 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1924
timestamp 1666464484
transform 1 0 49056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1925
timestamp 1666464484
transform 1 0 57008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1926
timestamp 1666464484
transform 1 0 64960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1927
timestamp 1666464484
transform 1 0 72912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1928
timestamp 1666464484
transform 1 0 80864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1929
timestamp 1666464484
transform 1 0 88816 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1930
timestamp 1666464484
transform 1 0 96768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1931
timestamp 1666464484
transform 1 0 104720 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1932
timestamp 1666464484
transform 1 0 112672 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1933
timestamp 1666464484
transform 1 0 120624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1934
timestamp 1666464484
transform 1 0 128576 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1935
timestamp 1666464484
transform 1 0 136528 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1936
timestamp 1666464484
transform 1 0 144480 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1937
timestamp 1666464484
transform 1 0 152432 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1938
timestamp 1666464484
transform 1 0 160384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1939
timestamp 1666464484
transform 1 0 168336 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1940
timestamp 1666464484
transform 1 0 176288 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1941
timestamp 1666464484
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1942
timestamp 1666464484
transform 1 0 13216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1943
timestamp 1666464484
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1944
timestamp 1666464484
transform 1 0 29120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1945
timestamp 1666464484
transform 1 0 37072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1946
timestamp 1666464484
transform 1 0 45024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1947
timestamp 1666464484
transform 1 0 52976 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1948
timestamp 1666464484
transform 1 0 60928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1949
timestamp 1666464484
transform 1 0 68880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1950
timestamp 1666464484
transform 1 0 76832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1951
timestamp 1666464484
transform 1 0 84784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1952
timestamp 1666464484
transform 1 0 92736 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1953
timestamp 1666464484
transform 1 0 100688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1954
timestamp 1666464484
transform 1 0 108640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1955
timestamp 1666464484
transform 1 0 116592 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1956
timestamp 1666464484
transform 1 0 124544 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1957
timestamp 1666464484
transform 1 0 132496 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1958
timestamp 1666464484
transform 1 0 140448 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1959
timestamp 1666464484
transform 1 0 148400 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1960
timestamp 1666464484
transform 1 0 156352 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1961
timestamp 1666464484
transform 1 0 164304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1962
timestamp 1666464484
transform 1 0 172256 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1963
timestamp 1666464484
transform 1 0 9296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1964
timestamp 1666464484
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1965
timestamp 1666464484
transform 1 0 25200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1966
timestamp 1666464484
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1967
timestamp 1666464484
transform 1 0 41104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1968
timestamp 1666464484
transform 1 0 49056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1969
timestamp 1666464484
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1970
timestamp 1666464484
transform 1 0 64960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1971
timestamp 1666464484
transform 1 0 72912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1972
timestamp 1666464484
transform 1 0 80864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1973
timestamp 1666464484
transform 1 0 88816 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1974
timestamp 1666464484
transform 1 0 96768 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1975
timestamp 1666464484
transform 1 0 104720 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1976
timestamp 1666464484
transform 1 0 112672 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1977
timestamp 1666464484
transform 1 0 120624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1978
timestamp 1666464484
transform 1 0 128576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1979
timestamp 1666464484
transform 1 0 136528 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1980
timestamp 1666464484
transform 1 0 144480 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1981
timestamp 1666464484
transform 1 0 152432 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1982
timestamp 1666464484
transform 1 0 160384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1983
timestamp 1666464484
transform 1 0 168336 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1984
timestamp 1666464484
transform 1 0 176288 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1985
timestamp 1666464484
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1986
timestamp 1666464484
transform 1 0 13216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1987
timestamp 1666464484
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1988
timestamp 1666464484
transform 1 0 29120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1989
timestamp 1666464484
transform 1 0 37072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1990
timestamp 1666464484
transform 1 0 45024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1991
timestamp 1666464484
transform 1 0 52976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1992
timestamp 1666464484
transform 1 0 60928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1993
timestamp 1666464484
transform 1 0 68880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1994
timestamp 1666464484
transform 1 0 76832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1995
timestamp 1666464484
transform 1 0 84784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1996
timestamp 1666464484
transform 1 0 92736 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1997
timestamp 1666464484
transform 1 0 100688 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1998
timestamp 1666464484
transform 1 0 108640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1999
timestamp 1666464484
transform 1 0 116592 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2000
timestamp 1666464484
transform 1 0 124544 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2001
timestamp 1666464484
transform 1 0 132496 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2002
timestamp 1666464484
transform 1 0 140448 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2003
timestamp 1666464484
transform 1 0 148400 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2004
timestamp 1666464484
transform 1 0 156352 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2005
timestamp 1666464484
transform 1 0 164304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2006
timestamp 1666464484
transform 1 0 172256 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2007
timestamp 1666464484
transform 1 0 9296 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2008
timestamp 1666464484
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2009
timestamp 1666464484
transform 1 0 25200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2010
timestamp 1666464484
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2011
timestamp 1666464484
transform 1 0 41104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2012
timestamp 1666464484
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2013
timestamp 1666464484
transform 1 0 57008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2014
timestamp 1666464484
transform 1 0 64960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2015
timestamp 1666464484
transform 1 0 72912 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2016
timestamp 1666464484
transform 1 0 80864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2017
timestamp 1666464484
transform 1 0 88816 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2018
timestamp 1666464484
transform 1 0 96768 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2019
timestamp 1666464484
transform 1 0 104720 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2020
timestamp 1666464484
transform 1 0 112672 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2021
timestamp 1666464484
transform 1 0 120624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2022
timestamp 1666464484
transform 1 0 128576 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2023
timestamp 1666464484
transform 1 0 136528 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2024
timestamp 1666464484
transform 1 0 144480 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2025
timestamp 1666464484
transform 1 0 152432 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2026
timestamp 1666464484
transform 1 0 160384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2027
timestamp 1666464484
transform 1 0 168336 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2028
timestamp 1666464484
transform 1 0 176288 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2029
timestamp 1666464484
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2030
timestamp 1666464484
transform 1 0 13216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2031
timestamp 1666464484
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2032
timestamp 1666464484
transform 1 0 29120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2033
timestamp 1666464484
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2034
timestamp 1666464484
transform 1 0 45024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2035
timestamp 1666464484
transform 1 0 52976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2036
timestamp 1666464484
transform 1 0 60928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2037
timestamp 1666464484
transform 1 0 68880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2038
timestamp 1666464484
transform 1 0 76832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2039
timestamp 1666464484
transform 1 0 84784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2040
timestamp 1666464484
transform 1 0 92736 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2041
timestamp 1666464484
transform 1 0 100688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2042
timestamp 1666464484
transform 1 0 108640 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2043
timestamp 1666464484
transform 1 0 116592 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2044
timestamp 1666464484
transform 1 0 124544 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2045
timestamp 1666464484
transform 1 0 132496 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2046
timestamp 1666464484
transform 1 0 140448 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2047
timestamp 1666464484
transform 1 0 148400 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2048
timestamp 1666464484
transform 1 0 156352 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2049
timestamp 1666464484
transform 1 0 164304 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2050
timestamp 1666464484
transform 1 0 172256 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2051
timestamp 1666464484
transform 1 0 9296 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2052
timestamp 1666464484
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2053
timestamp 1666464484
transform 1 0 25200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2054
timestamp 1666464484
transform 1 0 33152 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2055
timestamp 1666464484
transform 1 0 41104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2056
timestamp 1666464484
transform 1 0 49056 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2057
timestamp 1666464484
transform 1 0 57008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2058
timestamp 1666464484
transform 1 0 64960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2059
timestamp 1666464484
transform 1 0 72912 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2060
timestamp 1666464484
transform 1 0 80864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2061
timestamp 1666464484
transform 1 0 88816 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2062
timestamp 1666464484
transform 1 0 96768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2063
timestamp 1666464484
transform 1 0 104720 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2064
timestamp 1666464484
transform 1 0 112672 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2065
timestamp 1666464484
transform 1 0 120624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2066
timestamp 1666464484
transform 1 0 128576 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2067
timestamp 1666464484
transform 1 0 136528 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2068
timestamp 1666464484
transform 1 0 144480 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2069
timestamp 1666464484
transform 1 0 152432 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2070
timestamp 1666464484
transform 1 0 160384 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2071
timestamp 1666464484
transform 1 0 168336 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2072
timestamp 1666464484
transform 1 0 176288 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2073
timestamp 1666464484
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2074
timestamp 1666464484
transform 1 0 13216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2075
timestamp 1666464484
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2076
timestamp 1666464484
transform 1 0 29120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2077
timestamp 1666464484
transform 1 0 37072 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2078
timestamp 1666464484
transform 1 0 45024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2079
timestamp 1666464484
transform 1 0 52976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2080
timestamp 1666464484
transform 1 0 60928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2081
timestamp 1666464484
transform 1 0 68880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2082
timestamp 1666464484
transform 1 0 76832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2083
timestamp 1666464484
transform 1 0 84784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2084
timestamp 1666464484
transform 1 0 92736 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2085
timestamp 1666464484
transform 1 0 100688 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2086
timestamp 1666464484
transform 1 0 108640 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2087
timestamp 1666464484
transform 1 0 116592 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2088
timestamp 1666464484
transform 1 0 124544 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2089
timestamp 1666464484
transform 1 0 132496 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2090
timestamp 1666464484
transform 1 0 140448 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2091
timestamp 1666464484
transform 1 0 148400 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2092
timestamp 1666464484
transform 1 0 156352 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2093
timestamp 1666464484
transform 1 0 164304 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2094
timestamp 1666464484
transform 1 0 172256 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2095
timestamp 1666464484
transform 1 0 9296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2096
timestamp 1666464484
transform 1 0 17248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2097
timestamp 1666464484
transform 1 0 25200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2098
timestamp 1666464484
transform 1 0 33152 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2099
timestamp 1666464484
transform 1 0 41104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2100
timestamp 1666464484
transform 1 0 49056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2101
timestamp 1666464484
transform 1 0 57008 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2102
timestamp 1666464484
transform 1 0 64960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2103
timestamp 1666464484
transform 1 0 72912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2104
timestamp 1666464484
transform 1 0 80864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2105
timestamp 1666464484
transform 1 0 88816 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2106
timestamp 1666464484
transform 1 0 96768 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2107
timestamp 1666464484
transform 1 0 104720 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2108
timestamp 1666464484
transform 1 0 112672 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2109
timestamp 1666464484
transform 1 0 120624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2110
timestamp 1666464484
transform 1 0 128576 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2111
timestamp 1666464484
transform 1 0 136528 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2112
timestamp 1666464484
transform 1 0 144480 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2113
timestamp 1666464484
transform 1 0 152432 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2114
timestamp 1666464484
transform 1 0 160384 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2115
timestamp 1666464484
transform 1 0 168336 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2116
timestamp 1666464484
transform 1 0 176288 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2117
timestamp 1666464484
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2118
timestamp 1666464484
transform 1 0 13216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2119
timestamp 1666464484
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2120
timestamp 1666464484
transform 1 0 29120 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2121
timestamp 1666464484
transform 1 0 37072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2122
timestamp 1666464484
transform 1 0 45024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2123
timestamp 1666464484
transform 1 0 52976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2124
timestamp 1666464484
transform 1 0 60928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2125
timestamp 1666464484
transform 1 0 68880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2126
timestamp 1666464484
transform 1 0 76832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2127
timestamp 1666464484
transform 1 0 84784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2128
timestamp 1666464484
transform 1 0 92736 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2129
timestamp 1666464484
transform 1 0 100688 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2130
timestamp 1666464484
transform 1 0 108640 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2131
timestamp 1666464484
transform 1 0 116592 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2132
timestamp 1666464484
transform 1 0 124544 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2133
timestamp 1666464484
transform 1 0 132496 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2134
timestamp 1666464484
transform 1 0 140448 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2135
timestamp 1666464484
transform 1 0 148400 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2136
timestamp 1666464484
transform 1 0 156352 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2137
timestamp 1666464484
transform 1 0 164304 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2138
timestamp 1666464484
transform 1 0 172256 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2139
timestamp 1666464484
transform 1 0 9296 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2140
timestamp 1666464484
transform 1 0 17248 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2141
timestamp 1666464484
transform 1 0 25200 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2142
timestamp 1666464484
transform 1 0 33152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2143
timestamp 1666464484
transform 1 0 41104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2144
timestamp 1666464484
transform 1 0 49056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2145
timestamp 1666464484
transform 1 0 57008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2146
timestamp 1666464484
transform 1 0 64960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2147
timestamp 1666464484
transform 1 0 72912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2148
timestamp 1666464484
transform 1 0 80864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2149
timestamp 1666464484
transform 1 0 88816 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2150
timestamp 1666464484
transform 1 0 96768 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2151
timestamp 1666464484
transform 1 0 104720 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2152
timestamp 1666464484
transform 1 0 112672 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2153
timestamp 1666464484
transform 1 0 120624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2154
timestamp 1666464484
transform 1 0 128576 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2155
timestamp 1666464484
transform 1 0 136528 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2156
timestamp 1666464484
transform 1 0 144480 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2157
timestamp 1666464484
transform 1 0 152432 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2158
timestamp 1666464484
transform 1 0 160384 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2159
timestamp 1666464484
transform 1 0 168336 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2160
timestamp 1666464484
transform 1 0 176288 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2161
timestamp 1666464484
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2162
timestamp 1666464484
transform 1 0 13216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2163
timestamp 1666464484
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2164
timestamp 1666464484
transform 1 0 29120 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2165
timestamp 1666464484
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2166
timestamp 1666464484
transform 1 0 45024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2167
timestamp 1666464484
transform 1 0 52976 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2168
timestamp 1666464484
transform 1 0 60928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2169
timestamp 1666464484
transform 1 0 68880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2170
timestamp 1666464484
transform 1 0 76832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2171
timestamp 1666464484
transform 1 0 84784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2172
timestamp 1666464484
transform 1 0 92736 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2173
timestamp 1666464484
transform 1 0 100688 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2174
timestamp 1666464484
transform 1 0 108640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2175
timestamp 1666464484
transform 1 0 116592 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2176
timestamp 1666464484
transform 1 0 124544 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2177
timestamp 1666464484
transform 1 0 132496 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2178
timestamp 1666464484
transform 1 0 140448 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2179
timestamp 1666464484
transform 1 0 148400 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2180
timestamp 1666464484
transform 1 0 156352 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2181
timestamp 1666464484
transform 1 0 164304 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2182
timestamp 1666464484
transform 1 0 172256 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2183
timestamp 1666464484
transform 1 0 9296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2184
timestamp 1666464484
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2185
timestamp 1666464484
transform 1 0 25200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2186
timestamp 1666464484
transform 1 0 33152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2187
timestamp 1666464484
transform 1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2188
timestamp 1666464484
transform 1 0 49056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2189
timestamp 1666464484
transform 1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2190
timestamp 1666464484
transform 1 0 64960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2191
timestamp 1666464484
transform 1 0 72912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2192
timestamp 1666464484
transform 1 0 80864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2193
timestamp 1666464484
transform 1 0 88816 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2194
timestamp 1666464484
transform 1 0 96768 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2195
timestamp 1666464484
transform 1 0 104720 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2196
timestamp 1666464484
transform 1 0 112672 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2197
timestamp 1666464484
transform 1 0 120624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2198
timestamp 1666464484
transform 1 0 128576 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2199
timestamp 1666464484
transform 1 0 136528 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2200
timestamp 1666464484
transform 1 0 144480 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2201
timestamp 1666464484
transform 1 0 152432 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2202
timestamp 1666464484
transform 1 0 160384 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2203
timestamp 1666464484
transform 1 0 168336 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2204
timestamp 1666464484
transform 1 0 176288 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2205
timestamp 1666464484
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2206
timestamp 1666464484
transform 1 0 13216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2207
timestamp 1666464484
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2208
timestamp 1666464484
transform 1 0 29120 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2209
timestamp 1666464484
transform 1 0 37072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2210
timestamp 1666464484
transform 1 0 45024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2211
timestamp 1666464484
transform 1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2212
timestamp 1666464484
transform 1 0 60928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2213
timestamp 1666464484
transform 1 0 68880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2214
timestamp 1666464484
transform 1 0 76832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2215
timestamp 1666464484
transform 1 0 84784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2216
timestamp 1666464484
transform 1 0 92736 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2217
timestamp 1666464484
transform 1 0 100688 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2218
timestamp 1666464484
transform 1 0 108640 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2219
timestamp 1666464484
transform 1 0 116592 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2220
timestamp 1666464484
transform 1 0 124544 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2221
timestamp 1666464484
transform 1 0 132496 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2222
timestamp 1666464484
transform 1 0 140448 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2223
timestamp 1666464484
transform 1 0 148400 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2224
timestamp 1666464484
transform 1 0 156352 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2225
timestamp 1666464484
transform 1 0 164304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2226
timestamp 1666464484
transform 1 0 172256 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2227
timestamp 1666464484
transform 1 0 9296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2228
timestamp 1666464484
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2229
timestamp 1666464484
transform 1 0 25200 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2230
timestamp 1666464484
transform 1 0 33152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2231
timestamp 1666464484
transform 1 0 41104 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2232
timestamp 1666464484
transform 1 0 49056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2233
timestamp 1666464484
transform 1 0 57008 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2234
timestamp 1666464484
transform 1 0 64960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2235
timestamp 1666464484
transform 1 0 72912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2236
timestamp 1666464484
transform 1 0 80864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2237
timestamp 1666464484
transform 1 0 88816 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2238
timestamp 1666464484
transform 1 0 96768 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2239
timestamp 1666464484
transform 1 0 104720 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2240
timestamp 1666464484
transform 1 0 112672 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2241
timestamp 1666464484
transform 1 0 120624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2242
timestamp 1666464484
transform 1 0 128576 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2243
timestamp 1666464484
transform 1 0 136528 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2244
timestamp 1666464484
transform 1 0 144480 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2245
timestamp 1666464484
transform 1 0 152432 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2246
timestamp 1666464484
transform 1 0 160384 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2247
timestamp 1666464484
transform 1 0 168336 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2248
timestamp 1666464484
transform 1 0 176288 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2249
timestamp 1666464484
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2250
timestamp 1666464484
transform 1 0 13216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2251
timestamp 1666464484
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2252
timestamp 1666464484
transform 1 0 29120 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2253
timestamp 1666464484
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2254
timestamp 1666464484
transform 1 0 45024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2255
timestamp 1666464484
transform 1 0 52976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2256
timestamp 1666464484
transform 1 0 60928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2257
timestamp 1666464484
transform 1 0 68880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2258
timestamp 1666464484
transform 1 0 76832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2259
timestamp 1666464484
transform 1 0 84784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2260
timestamp 1666464484
transform 1 0 92736 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2261
timestamp 1666464484
transform 1 0 100688 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2262
timestamp 1666464484
transform 1 0 108640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2263
timestamp 1666464484
transform 1 0 116592 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2264
timestamp 1666464484
transform 1 0 124544 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2265
timestamp 1666464484
transform 1 0 132496 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2266
timestamp 1666464484
transform 1 0 140448 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2267
timestamp 1666464484
transform 1 0 148400 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2268
timestamp 1666464484
transform 1 0 156352 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2269
timestamp 1666464484
transform 1 0 164304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2270
timestamp 1666464484
transform 1 0 172256 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2271
timestamp 1666464484
transform 1 0 9296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2272
timestamp 1666464484
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2273
timestamp 1666464484
transform 1 0 25200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2274
timestamp 1666464484
transform 1 0 33152 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2275
timestamp 1666464484
transform 1 0 41104 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2276
timestamp 1666464484
transform 1 0 49056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2277
timestamp 1666464484
transform 1 0 57008 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2278
timestamp 1666464484
transform 1 0 64960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2279
timestamp 1666464484
transform 1 0 72912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2280
timestamp 1666464484
transform 1 0 80864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2281
timestamp 1666464484
transform 1 0 88816 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2282
timestamp 1666464484
transform 1 0 96768 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2283
timestamp 1666464484
transform 1 0 104720 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2284
timestamp 1666464484
transform 1 0 112672 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2285
timestamp 1666464484
transform 1 0 120624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2286
timestamp 1666464484
transform 1 0 128576 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2287
timestamp 1666464484
transform 1 0 136528 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2288
timestamp 1666464484
transform 1 0 144480 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2289
timestamp 1666464484
transform 1 0 152432 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2290
timestamp 1666464484
transform 1 0 160384 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2291
timestamp 1666464484
transform 1 0 168336 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2292
timestamp 1666464484
transform 1 0 176288 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2293
timestamp 1666464484
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2294
timestamp 1666464484
transform 1 0 13216 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2295
timestamp 1666464484
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2296
timestamp 1666464484
transform 1 0 29120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2297
timestamp 1666464484
transform 1 0 37072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2298
timestamp 1666464484
transform 1 0 45024 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2299
timestamp 1666464484
transform 1 0 52976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2300
timestamp 1666464484
transform 1 0 60928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2301
timestamp 1666464484
transform 1 0 68880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2302
timestamp 1666464484
transform 1 0 76832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2303
timestamp 1666464484
transform 1 0 84784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2304
timestamp 1666464484
transform 1 0 92736 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2305
timestamp 1666464484
transform 1 0 100688 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2306
timestamp 1666464484
transform 1 0 108640 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2307
timestamp 1666464484
transform 1 0 116592 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2308
timestamp 1666464484
transform 1 0 124544 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2309
timestamp 1666464484
transform 1 0 132496 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2310
timestamp 1666464484
transform 1 0 140448 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2311
timestamp 1666464484
transform 1 0 148400 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2312
timestamp 1666464484
transform 1 0 156352 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2313
timestamp 1666464484
transform 1 0 164304 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2314
timestamp 1666464484
transform 1 0 172256 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2315
timestamp 1666464484
transform 1 0 9296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2316
timestamp 1666464484
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2317
timestamp 1666464484
transform 1 0 25200 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2318
timestamp 1666464484
transform 1 0 33152 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2319
timestamp 1666464484
transform 1 0 41104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2320
timestamp 1666464484
transform 1 0 49056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2321
timestamp 1666464484
transform 1 0 57008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2322
timestamp 1666464484
transform 1 0 64960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2323
timestamp 1666464484
transform 1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2324
timestamp 1666464484
transform 1 0 80864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2325
timestamp 1666464484
transform 1 0 88816 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2326
timestamp 1666464484
transform 1 0 96768 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2327
timestamp 1666464484
transform 1 0 104720 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2328
timestamp 1666464484
transform 1 0 112672 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2329
timestamp 1666464484
transform 1 0 120624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2330
timestamp 1666464484
transform 1 0 128576 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2331
timestamp 1666464484
transform 1 0 136528 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2332
timestamp 1666464484
transform 1 0 144480 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2333
timestamp 1666464484
transform 1 0 152432 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2334
timestamp 1666464484
transform 1 0 160384 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2335
timestamp 1666464484
transform 1 0 168336 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2336
timestamp 1666464484
transform 1 0 176288 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2337
timestamp 1666464484
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2338
timestamp 1666464484
transform 1 0 13216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2339
timestamp 1666464484
transform 1 0 21168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2340
timestamp 1666464484
transform 1 0 29120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2341
timestamp 1666464484
transform 1 0 37072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2342
timestamp 1666464484
transform 1 0 45024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2343
timestamp 1666464484
transform 1 0 52976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2344
timestamp 1666464484
transform 1 0 60928 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2345
timestamp 1666464484
transform 1 0 68880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2346
timestamp 1666464484
transform 1 0 76832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2347
timestamp 1666464484
transform 1 0 84784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2348
timestamp 1666464484
transform 1 0 92736 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2349
timestamp 1666464484
transform 1 0 100688 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2350
timestamp 1666464484
transform 1 0 108640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2351
timestamp 1666464484
transform 1 0 116592 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2352
timestamp 1666464484
transform 1 0 124544 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2353
timestamp 1666464484
transform 1 0 132496 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2354
timestamp 1666464484
transform 1 0 140448 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2355
timestamp 1666464484
transform 1 0 148400 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2356
timestamp 1666464484
transform 1 0 156352 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2357
timestamp 1666464484
transform 1 0 164304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2358
timestamp 1666464484
transform 1 0 172256 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2359
timestamp 1666464484
transform 1 0 9296 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2360
timestamp 1666464484
transform 1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2361
timestamp 1666464484
transform 1 0 25200 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2362
timestamp 1666464484
transform 1 0 33152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2363
timestamp 1666464484
transform 1 0 41104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2364
timestamp 1666464484
transform 1 0 49056 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2365
timestamp 1666464484
transform 1 0 57008 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2366
timestamp 1666464484
transform 1 0 64960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2367
timestamp 1666464484
transform 1 0 72912 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2368
timestamp 1666464484
transform 1 0 80864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2369
timestamp 1666464484
transform 1 0 88816 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2370
timestamp 1666464484
transform 1 0 96768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2371
timestamp 1666464484
transform 1 0 104720 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2372
timestamp 1666464484
transform 1 0 112672 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2373
timestamp 1666464484
transform 1 0 120624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2374
timestamp 1666464484
transform 1 0 128576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2375
timestamp 1666464484
transform 1 0 136528 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2376
timestamp 1666464484
transform 1 0 144480 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2377
timestamp 1666464484
transform 1 0 152432 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2378
timestamp 1666464484
transform 1 0 160384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2379
timestamp 1666464484
transform 1 0 168336 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2380
timestamp 1666464484
transform 1 0 176288 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2381
timestamp 1666464484
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2382
timestamp 1666464484
transform 1 0 13216 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2383
timestamp 1666464484
transform 1 0 21168 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2384
timestamp 1666464484
transform 1 0 29120 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2385
timestamp 1666464484
transform 1 0 37072 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2386
timestamp 1666464484
transform 1 0 45024 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2387
timestamp 1666464484
transform 1 0 52976 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2388
timestamp 1666464484
transform 1 0 60928 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2389
timestamp 1666464484
transform 1 0 68880 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2390
timestamp 1666464484
transform 1 0 76832 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2391
timestamp 1666464484
transform 1 0 84784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2392
timestamp 1666464484
transform 1 0 92736 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2393
timestamp 1666464484
transform 1 0 100688 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2394
timestamp 1666464484
transform 1 0 108640 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2395
timestamp 1666464484
transform 1 0 116592 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2396
timestamp 1666464484
transform 1 0 124544 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2397
timestamp 1666464484
transform 1 0 132496 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2398
timestamp 1666464484
transform 1 0 140448 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2399
timestamp 1666464484
transform 1 0 148400 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2400
timestamp 1666464484
transform 1 0 156352 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2401
timestamp 1666464484
transform 1 0 164304 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2402
timestamp 1666464484
transform 1 0 172256 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2403
timestamp 1666464484
transform 1 0 9296 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2404
timestamp 1666464484
transform 1 0 17248 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2405
timestamp 1666464484
transform 1 0 25200 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2406
timestamp 1666464484
transform 1 0 33152 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2407
timestamp 1666464484
transform 1 0 41104 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2408
timestamp 1666464484
transform 1 0 49056 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2409
timestamp 1666464484
transform 1 0 57008 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2410
timestamp 1666464484
transform 1 0 64960 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2411
timestamp 1666464484
transform 1 0 72912 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2412
timestamp 1666464484
transform 1 0 80864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2413
timestamp 1666464484
transform 1 0 88816 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2414
timestamp 1666464484
transform 1 0 96768 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2415
timestamp 1666464484
transform 1 0 104720 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2416
timestamp 1666464484
transform 1 0 112672 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2417
timestamp 1666464484
transform 1 0 120624 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2418
timestamp 1666464484
transform 1 0 128576 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2419
timestamp 1666464484
transform 1 0 136528 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2420
timestamp 1666464484
transform 1 0 144480 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2421
timestamp 1666464484
transform 1 0 152432 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2422
timestamp 1666464484
transform 1 0 160384 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2423
timestamp 1666464484
transform 1 0 168336 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2424
timestamp 1666464484
transform 1 0 176288 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2425
timestamp 1666464484
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2426
timestamp 1666464484
transform 1 0 13216 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2427
timestamp 1666464484
transform 1 0 21168 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2428
timestamp 1666464484
transform 1 0 29120 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2429
timestamp 1666464484
transform 1 0 37072 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2430
timestamp 1666464484
transform 1 0 45024 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2431
timestamp 1666464484
transform 1 0 52976 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2432
timestamp 1666464484
transform 1 0 60928 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2433
timestamp 1666464484
transform 1 0 68880 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2434
timestamp 1666464484
transform 1 0 76832 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2435
timestamp 1666464484
transform 1 0 84784 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2436
timestamp 1666464484
transform 1 0 92736 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2437
timestamp 1666464484
transform 1 0 100688 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2438
timestamp 1666464484
transform 1 0 108640 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2439
timestamp 1666464484
transform 1 0 116592 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2440
timestamp 1666464484
transform 1 0 124544 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2441
timestamp 1666464484
transform 1 0 132496 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2442
timestamp 1666464484
transform 1 0 140448 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2443
timestamp 1666464484
transform 1 0 148400 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2444
timestamp 1666464484
transform 1 0 156352 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2445
timestamp 1666464484
transform 1 0 164304 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2446
timestamp 1666464484
transform 1 0 172256 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2447
timestamp 1666464484
transform 1 0 9296 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2448
timestamp 1666464484
transform 1 0 17248 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2449
timestamp 1666464484
transform 1 0 25200 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2450
timestamp 1666464484
transform 1 0 33152 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2451
timestamp 1666464484
transform 1 0 41104 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2452
timestamp 1666464484
transform 1 0 49056 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2453
timestamp 1666464484
transform 1 0 57008 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2454
timestamp 1666464484
transform 1 0 64960 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2455
timestamp 1666464484
transform 1 0 72912 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2456
timestamp 1666464484
transform 1 0 80864 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2457
timestamp 1666464484
transform 1 0 88816 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2458
timestamp 1666464484
transform 1 0 96768 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2459
timestamp 1666464484
transform 1 0 104720 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2460
timestamp 1666464484
transform 1 0 112672 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2461
timestamp 1666464484
transform 1 0 120624 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2462
timestamp 1666464484
transform 1 0 128576 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2463
timestamp 1666464484
transform 1 0 136528 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2464
timestamp 1666464484
transform 1 0 144480 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2465
timestamp 1666464484
transform 1 0 152432 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2466
timestamp 1666464484
transform 1 0 160384 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2467
timestamp 1666464484
transform 1 0 168336 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2468
timestamp 1666464484
transform 1 0 176288 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2469
timestamp 1666464484
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2470
timestamp 1666464484
transform 1 0 13216 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2471
timestamp 1666464484
transform 1 0 21168 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2472
timestamp 1666464484
transform 1 0 29120 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2473
timestamp 1666464484
transform 1 0 37072 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2474
timestamp 1666464484
transform 1 0 45024 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2475
timestamp 1666464484
transform 1 0 52976 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2476
timestamp 1666464484
transform 1 0 60928 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2477
timestamp 1666464484
transform 1 0 68880 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2478
timestamp 1666464484
transform 1 0 76832 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2479
timestamp 1666464484
transform 1 0 84784 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2480
timestamp 1666464484
transform 1 0 92736 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2481
timestamp 1666464484
transform 1 0 100688 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2482
timestamp 1666464484
transform 1 0 108640 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2483
timestamp 1666464484
transform 1 0 116592 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2484
timestamp 1666464484
transform 1 0 124544 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2485
timestamp 1666464484
transform 1 0 132496 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2486
timestamp 1666464484
transform 1 0 140448 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2487
timestamp 1666464484
transform 1 0 148400 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2488
timestamp 1666464484
transform 1 0 156352 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2489
timestamp 1666464484
transform 1 0 164304 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2490
timestamp 1666464484
transform 1 0 172256 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2491
timestamp 1666464484
transform 1 0 9296 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2492
timestamp 1666464484
transform 1 0 17248 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2493
timestamp 1666464484
transform 1 0 25200 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2494
timestamp 1666464484
transform 1 0 33152 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2495
timestamp 1666464484
transform 1 0 41104 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2496
timestamp 1666464484
transform 1 0 49056 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2497
timestamp 1666464484
transform 1 0 57008 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2498
timestamp 1666464484
transform 1 0 64960 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2499
timestamp 1666464484
transform 1 0 72912 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2500
timestamp 1666464484
transform 1 0 80864 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2501
timestamp 1666464484
transform 1 0 88816 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2502
timestamp 1666464484
transform 1 0 96768 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2503
timestamp 1666464484
transform 1 0 104720 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2504
timestamp 1666464484
transform 1 0 112672 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2505
timestamp 1666464484
transform 1 0 120624 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2506
timestamp 1666464484
transform 1 0 128576 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2507
timestamp 1666464484
transform 1 0 136528 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2508
timestamp 1666464484
transform 1 0 144480 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2509
timestamp 1666464484
transform 1 0 152432 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2510
timestamp 1666464484
transform 1 0 160384 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2511
timestamp 1666464484
transform 1 0 168336 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2512
timestamp 1666464484
transform 1 0 176288 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2513
timestamp 1666464484
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2514
timestamp 1666464484
transform 1 0 13216 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2515
timestamp 1666464484
transform 1 0 21168 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2516
timestamp 1666464484
transform 1 0 29120 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2517
timestamp 1666464484
transform 1 0 37072 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2518
timestamp 1666464484
transform 1 0 45024 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2519
timestamp 1666464484
transform 1 0 52976 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2520
timestamp 1666464484
transform 1 0 60928 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2521
timestamp 1666464484
transform 1 0 68880 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2522
timestamp 1666464484
transform 1 0 76832 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2523
timestamp 1666464484
transform 1 0 84784 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2524
timestamp 1666464484
transform 1 0 92736 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2525
timestamp 1666464484
transform 1 0 100688 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2526
timestamp 1666464484
transform 1 0 108640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2527
timestamp 1666464484
transform 1 0 116592 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2528
timestamp 1666464484
transform 1 0 124544 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2529
timestamp 1666464484
transform 1 0 132496 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2530
timestamp 1666464484
transform 1 0 140448 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2531
timestamp 1666464484
transform 1 0 148400 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2532
timestamp 1666464484
transform 1 0 156352 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2533
timestamp 1666464484
transform 1 0 164304 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2534
timestamp 1666464484
transform 1 0 172256 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2535
timestamp 1666464484
transform 1 0 9296 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2536
timestamp 1666464484
transform 1 0 17248 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2537
timestamp 1666464484
transform 1 0 25200 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2538
timestamp 1666464484
transform 1 0 33152 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2539
timestamp 1666464484
transform 1 0 41104 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2540
timestamp 1666464484
transform 1 0 49056 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2541
timestamp 1666464484
transform 1 0 57008 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2542
timestamp 1666464484
transform 1 0 64960 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2543
timestamp 1666464484
transform 1 0 72912 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2544
timestamp 1666464484
transform 1 0 80864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2545
timestamp 1666464484
transform 1 0 88816 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2546
timestamp 1666464484
transform 1 0 96768 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2547
timestamp 1666464484
transform 1 0 104720 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2548
timestamp 1666464484
transform 1 0 112672 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2549
timestamp 1666464484
transform 1 0 120624 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2550
timestamp 1666464484
transform 1 0 128576 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2551
timestamp 1666464484
transform 1 0 136528 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2552
timestamp 1666464484
transform 1 0 144480 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2553
timestamp 1666464484
transform 1 0 152432 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2554
timestamp 1666464484
transform 1 0 160384 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2555
timestamp 1666464484
transform 1 0 168336 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2556
timestamp 1666464484
transform 1 0 176288 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2557
timestamp 1666464484
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2558
timestamp 1666464484
transform 1 0 13216 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2559
timestamp 1666464484
transform 1 0 21168 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2560
timestamp 1666464484
transform 1 0 29120 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2561
timestamp 1666464484
transform 1 0 37072 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2562
timestamp 1666464484
transform 1 0 45024 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2563
timestamp 1666464484
transform 1 0 52976 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2564
timestamp 1666464484
transform 1 0 60928 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2565
timestamp 1666464484
transform 1 0 68880 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2566
timestamp 1666464484
transform 1 0 76832 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2567
timestamp 1666464484
transform 1 0 84784 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2568
timestamp 1666464484
transform 1 0 92736 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2569
timestamp 1666464484
transform 1 0 100688 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2570
timestamp 1666464484
transform 1 0 108640 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2571
timestamp 1666464484
transform 1 0 116592 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2572
timestamp 1666464484
transform 1 0 124544 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2573
timestamp 1666464484
transform 1 0 132496 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2574
timestamp 1666464484
transform 1 0 140448 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2575
timestamp 1666464484
transform 1 0 148400 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2576
timestamp 1666464484
transform 1 0 156352 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2577
timestamp 1666464484
transform 1 0 164304 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2578
timestamp 1666464484
transform 1 0 172256 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2579
timestamp 1666464484
transform 1 0 9296 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2580
timestamp 1666464484
transform 1 0 17248 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2581
timestamp 1666464484
transform 1 0 25200 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2582
timestamp 1666464484
transform 1 0 33152 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2583
timestamp 1666464484
transform 1 0 41104 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2584
timestamp 1666464484
transform 1 0 49056 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2585
timestamp 1666464484
transform 1 0 57008 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2586
timestamp 1666464484
transform 1 0 64960 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2587
timestamp 1666464484
transform 1 0 72912 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2588
timestamp 1666464484
transform 1 0 80864 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2589
timestamp 1666464484
transform 1 0 88816 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2590
timestamp 1666464484
transform 1 0 96768 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2591
timestamp 1666464484
transform 1 0 104720 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2592
timestamp 1666464484
transform 1 0 112672 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2593
timestamp 1666464484
transform 1 0 120624 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2594
timestamp 1666464484
transform 1 0 128576 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2595
timestamp 1666464484
transform 1 0 136528 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2596
timestamp 1666464484
transform 1 0 144480 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2597
timestamp 1666464484
transform 1 0 152432 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2598
timestamp 1666464484
transform 1 0 160384 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2599
timestamp 1666464484
transform 1 0 168336 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2600
timestamp 1666464484
transform 1 0 176288 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2601
timestamp 1666464484
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2602
timestamp 1666464484
transform 1 0 13216 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2603
timestamp 1666464484
transform 1 0 21168 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2604
timestamp 1666464484
transform 1 0 29120 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2605
timestamp 1666464484
transform 1 0 37072 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2606
timestamp 1666464484
transform 1 0 45024 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2607
timestamp 1666464484
transform 1 0 52976 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2608
timestamp 1666464484
transform 1 0 60928 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2609
timestamp 1666464484
transform 1 0 68880 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2610
timestamp 1666464484
transform 1 0 76832 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2611
timestamp 1666464484
transform 1 0 84784 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2612
timestamp 1666464484
transform 1 0 92736 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2613
timestamp 1666464484
transform 1 0 100688 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2614
timestamp 1666464484
transform 1 0 108640 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2615
timestamp 1666464484
transform 1 0 116592 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2616
timestamp 1666464484
transform 1 0 124544 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2617
timestamp 1666464484
transform 1 0 132496 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2618
timestamp 1666464484
transform 1 0 140448 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2619
timestamp 1666464484
transform 1 0 148400 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2620
timestamp 1666464484
transform 1 0 156352 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2621
timestamp 1666464484
transform 1 0 164304 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2622
timestamp 1666464484
transform 1 0 172256 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2623
timestamp 1666464484
transform 1 0 9296 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2624
timestamp 1666464484
transform 1 0 17248 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2625
timestamp 1666464484
transform 1 0 25200 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2626
timestamp 1666464484
transform 1 0 33152 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2627
timestamp 1666464484
transform 1 0 41104 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2628
timestamp 1666464484
transform 1 0 49056 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2629
timestamp 1666464484
transform 1 0 57008 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2630
timestamp 1666464484
transform 1 0 64960 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2631
timestamp 1666464484
transform 1 0 72912 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2632
timestamp 1666464484
transform 1 0 80864 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2633
timestamp 1666464484
transform 1 0 88816 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2634
timestamp 1666464484
transform 1 0 96768 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2635
timestamp 1666464484
transform 1 0 104720 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2636
timestamp 1666464484
transform 1 0 112672 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2637
timestamp 1666464484
transform 1 0 120624 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2638
timestamp 1666464484
transform 1 0 128576 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2639
timestamp 1666464484
transform 1 0 136528 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2640
timestamp 1666464484
transform 1 0 144480 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2641
timestamp 1666464484
transform 1 0 152432 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2642
timestamp 1666464484
transform 1 0 160384 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2643
timestamp 1666464484
transform 1 0 168336 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2644
timestamp 1666464484
transform 1 0 176288 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2645
timestamp 1666464484
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2646
timestamp 1666464484
transform 1 0 13216 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2647
timestamp 1666464484
transform 1 0 21168 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2648
timestamp 1666464484
transform 1 0 29120 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2649
timestamp 1666464484
transform 1 0 37072 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2650
timestamp 1666464484
transform 1 0 45024 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2651
timestamp 1666464484
transform 1 0 52976 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2652
timestamp 1666464484
transform 1 0 60928 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2653
timestamp 1666464484
transform 1 0 68880 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2654
timestamp 1666464484
transform 1 0 76832 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2655
timestamp 1666464484
transform 1 0 84784 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2656
timestamp 1666464484
transform 1 0 92736 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2657
timestamp 1666464484
transform 1 0 100688 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2658
timestamp 1666464484
transform 1 0 108640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2659
timestamp 1666464484
transform 1 0 116592 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2660
timestamp 1666464484
transform 1 0 124544 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2661
timestamp 1666464484
transform 1 0 132496 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2662
timestamp 1666464484
transform 1 0 140448 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2663
timestamp 1666464484
transform 1 0 148400 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2664
timestamp 1666464484
transform 1 0 156352 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2665
timestamp 1666464484
transform 1 0 164304 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2666
timestamp 1666464484
transform 1 0 172256 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2667
timestamp 1666464484
transform 1 0 9296 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2668
timestamp 1666464484
transform 1 0 17248 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2669
timestamp 1666464484
transform 1 0 25200 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2670
timestamp 1666464484
transform 1 0 33152 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2671
timestamp 1666464484
transform 1 0 41104 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2672
timestamp 1666464484
transform 1 0 49056 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2673
timestamp 1666464484
transform 1 0 57008 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2674
timestamp 1666464484
transform 1 0 64960 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2675
timestamp 1666464484
transform 1 0 72912 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2676
timestamp 1666464484
transform 1 0 80864 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2677
timestamp 1666464484
transform 1 0 88816 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2678
timestamp 1666464484
transform 1 0 96768 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2679
timestamp 1666464484
transform 1 0 104720 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2680
timestamp 1666464484
transform 1 0 112672 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2681
timestamp 1666464484
transform 1 0 120624 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2682
timestamp 1666464484
transform 1 0 128576 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2683
timestamp 1666464484
transform 1 0 136528 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2684
timestamp 1666464484
transform 1 0 144480 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2685
timestamp 1666464484
transform 1 0 152432 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2686
timestamp 1666464484
transform 1 0 160384 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2687
timestamp 1666464484
transform 1 0 168336 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2688
timestamp 1666464484
transform 1 0 176288 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2689
timestamp 1666464484
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2690
timestamp 1666464484
transform 1 0 13216 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2691
timestamp 1666464484
transform 1 0 21168 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2692
timestamp 1666464484
transform 1 0 29120 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2693
timestamp 1666464484
transform 1 0 37072 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2694
timestamp 1666464484
transform 1 0 45024 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2695
timestamp 1666464484
transform 1 0 52976 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2696
timestamp 1666464484
transform 1 0 60928 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2697
timestamp 1666464484
transform 1 0 68880 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2698
timestamp 1666464484
transform 1 0 76832 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2699
timestamp 1666464484
transform 1 0 84784 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2700
timestamp 1666464484
transform 1 0 92736 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2701
timestamp 1666464484
transform 1 0 100688 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2702
timestamp 1666464484
transform 1 0 108640 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2703
timestamp 1666464484
transform 1 0 116592 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2704
timestamp 1666464484
transform 1 0 124544 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2705
timestamp 1666464484
transform 1 0 132496 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2706
timestamp 1666464484
transform 1 0 140448 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2707
timestamp 1666464484
transform 1 0 148400 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2708
timestamp 1666464484
transform 1 0 156352 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2709
timestamp 1666464484
transform 1 0 164304 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2710
timestamp 1666464484
transform 1 0 172256 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2711
timestamp 1666464484
transform 1 0 9296 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2712
timestamp 1666464484
transform 1 0 17248 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2713
timestamp 1666464484
transform 1 0 25200 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2714
timestamp 1666464484
transform 1 0 33152 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2715
timestamp 1666464484
transform 1 0 41104 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2716
timestamp 1666464484
transform 1 0 49056 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2717
timestamp 1666464484
transform 1 0 57008 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2718
timestamp 1666464484
transform 1 0 64960 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2719
timestamp 1666464484
transform 1 0 72912 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2720
timestamp 1666464484
transform 1 0 80864 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2721
timestamp 1666464484
transform 1 0 88816 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2722
timestamp 1666464484
transform 1 0 96768 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2723
timestamp 1666464484
transform 1 0 104720 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2724
timestamp 1666464484
transform 1 0 112672 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2725
timestamp 1666464484
transform 1 0 120624 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2726
timestamp 1666464484
transform 1 0 128576 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2727
timestamp 1666464484
transform 1 0 136528 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2728
timestamp 1666464484
transform 1 0 144480 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2729
timestamp 1666464484
transform 1 0 152432 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2730
timestamp 1666464484
transform 1 0 160384 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2731
timestamp 1666464484
transform 1 0 168336 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2732
timestamp 1666464484
transform 1 0 176288 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2733
timestamp 1666464484
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2734
timestamp 1666464484
transform 1 0 13216 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2735
timestamp 1666464484
transform 1 0 21168 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2736
timestamp 1666464484
transform 1 0 29120 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2737
timestamp 1666464484
transform 1 0 37072 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2738
timestamp 1666464484
transform 1 0 45024 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2739
timestamp 1666464484
transform 1 0 52976 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2740
timestamp 1666464484
transform 1 0 60928 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2741
timestamp 1666464484
transform 1 0 68880 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2742
timestamp 1666464484
transform 1 0 76832 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2743
timestamp 1666464484
transform 1 0 84784 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2744
timestamp 1666464484
transform 1 0 92736 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2745
timestamp 1666464484
transform 1 0 100688 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2746
timestamp 1666464484
transform 1 0 108640 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2747
timestamp 1666464484
transform 1 0 116592 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2748
timestamp 1666464484
transform 1 0 124544 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2749
timestamp 1666464484
transform 1 0 132496 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2750
timestamp 1666464484
transform 1 0 140448 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2751
timestamp 1666464484
transform 1 0 148400 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2752
timestamp 1666464484
transform 1 0 156352 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2753
timestamp 1666464484
transform 1 0 164304 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2754
timestamp 1666464484
transform 1 0 172256 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2755
timestamp 1666464484
transform 1 0 9296 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2756
timestamp 1666464484
transform 1 0 17248 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2757
timestamp 1666464484
transform 1 0 25200 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2758
timestamp 1666464484
transform 1 0 33152 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2759
timestamp 1666464484
transform 1 0 41104 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2760
timestamp 1666464484
transform 1 0 49056 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2761
timestamp 1666464484
transform 1 0 57008 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2762
timestamp 1666464484
transform 1 0 64960 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2763
timestamp 1666464484
transform 1 0 72912 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2764
timestamp 1666464484
transform 1 0 80864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2765
timestamp 1666464484
transform 1 0 88816 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2766
timestamp 1666464484
transform 1 0 96768 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2767
timestamp 1666464484
transform 1 0 104720 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2768
timestamp 1666464484
transform 1 0 112672 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2769
timestamp 1666464484
transform 1 0 120624 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2770
timestamp 1666464484
transform 1 0 128576 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2771
timestamp 1666464484
transform 1 0 136528 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2772
timestamp 1666464484
transform 1 0 144480 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2773
timestamp 1666464484
transform 1 0 152432 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2774
timestamp 1666464484
transform 1 0 160384 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2775
timestamp 1666464484
transform 1 0 168336 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2776
timestamp 1666464484
transform 1 0 176288 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2777
timestamp 1666464484
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2778
timestamp 1666464484
transform 1 0 13216 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2779
timestamp 1666464484
transform 1 0 21168 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2780
timestamp 1666464484
transform 1 0 29120 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2781
timestamp 1666464484
transform 1 0 37072 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2782
timestamp 1666464484
transform 1 0 45024 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2783
timestamp 1666464484
transform 1 0 52976 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2784
timestamp 1666464484
transform 1 0 60928 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2785
timestamp 1666464484
transform 1 0 68880 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2786
timestamp 1666464484
transform 1 0 76832 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2787
timestamp 1666464484
transform 1 0 84784 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2788
timestamp 1666464484
transform 1 0 92736 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2789
timestamp 1666464484
transform 1 0 100688 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2790
timestamp 1666464484
transform 1 0 108640 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2791
timestamp 1666464484
transform 1 0 116592 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2792
timestamp 1666464484
transform 1 0 124544 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2793
timestamp 1666464484
transform 1 0 132496 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2794
timestamp 1666464484
transform 1 0 140448 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2795
timestamp 1666464484
transform 1 0 148400 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2796
timestamp 1666464484
transform 1 0 156352 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2797
timestamp 1666464484
transform 1 0 164304 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2798
timestamp 1666464484
transform 1 0 172256 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2799
timestamp 1666464484
transform 1 0 9296 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2800
timestamp 1666464484
transform 1 0 17248 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2801
timestamp 1666464484
transform 1 0 25200 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2802
timestamp 1666464484
transform 1 0 33152 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2803
timestamp 1666464484
transform 1 0 41104 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2804
timestamp 1666464484
transform 1 0 49056 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2805
timestamp 1666464484
transform 1 0 57008 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2806
timestamp 1666464484
transform 1 0 64960 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2807
timestamp 1666464484
transform 1 0 72912 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2808
timestamp 1666464484
transform 1 0 80864 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2809
timestamp 1666464484
transform 1 0 88816 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2810
timestamp 1666464484
transform 1 0 96768 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2811
timestamp 1666464484
transform 1 0 104720 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2812
timestamp 1666464484
transform 1 0 112672 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2813
timestamp 1666464484
transform 1 0 120624 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2814
timestamp 1666464484
transform 1 0 128576 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2815
timestamp 1666464484
transform 1 0 136528 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2816
timestamp 1666464484
transform 1 0 144480 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2817
timestamp 1666464484
transform 1 0 152432 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2818
timestamp 1666464484
transform 1 0 160384 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2819
timestamp 1666464484
transform 1 0 168336 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2820
timestamp 1666464484
transform 1 0 176288 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2821
timestamp 1666464484
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2822
timestamp 1666464484
transform 1 0 13216 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2823
timestamp 1666464484
transform 1 0 21168 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2824
timestamp 1666464484
transform 1 0 29120 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2825
timestamp 1666464484
transform 1 0 37072 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2826
timestamp 1666464484
transform 1 0 45024 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2827
timestamp 1666464484
transform 1 0 52976 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2828
timestamp 1666464484
transform 1 0 60928 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2829
timestamp 1666464484
transform 1 0 68880 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2830
timestamp 1666464484
transform 1 0 76832 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2831
timestamp 1666464484
transform 1 0 84784 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2832
timestamp 1666464484
transform 1 0 92736 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2833
timestamp 1666464484
transform 1 0 100688 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2834
timestamp 1666464484
transform 1 0 108640 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2835
timestamp 1666464484
transform 1 0 116592 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2836
timestamp 1666464484
transform 1 0 124544 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2837
timestamp 1666464484
transform 1 0 132496 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2838
timestamp 1666464484
transform 1 0 140448 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2839
timestamp 1666464484
transform 1 0 148400 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2840
timestamp 1666464484
transform 1 0 156352 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2841
timestamp 1666464484
transform 1 0 164304 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2842
timestamp 1666464484
transform 1 0 172256 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2843
timestamp 1666464484
transform 1 0 9296 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2844
timestamp 1666464484
transform 1 0 17248 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2845
timestamp 1666464484
transform 1 0 25200 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2846
timestamp 1666464484
transform 1 0 33152 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2847
timestamp 1666464484
transform 1 0 41104 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2848
timestamp 1666464484
transform 1 0 49056 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2849
timestamp 1666464484
transform 1 0 57008 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2850
timestamp 1666464484
transform 1 0 64960 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2851
timestamp 1666464484
transform 1 0 72912 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2852
timestamp 1666464484
transform 1 0 80864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2853
timestamp 1666464484
transform 1 0 88816 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2854
timestamp 1666464484
transform 1 0 96768 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2855
timestamp 1666464484
transform 1 0 104720 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2856
timestamp 1666464484
transform 1 0 112672 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2857
timestamp 1666464484
transform 1 0 120624 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2858
timestamp 1666464484
transform 1 0 128576 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2859
timestamp 1666464484
transform 1 0 136528 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2860
timestamp 1666464484
transform 1 0 144480 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2861
timestamp 1666464484
transform 1 0 152432 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2862
timestamp 1666464484
transform 1 0 160384 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2863
timestamp 1666464484
transform 1 0 168336 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2864
timestamp 1666464484
transform 1 0 176288 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2865
timestamp 1666464484
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2866
timestamp 1666464484
transform 1 0 13216 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2867
timestamp 1666464484
transform 1 0 21168 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2868
timestamp 1666464484
transform 1 0 29120 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2869
timestamp 1666464484
transform 1 0 37072 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2870
timestamp 1666464484
transform 1 0 45024 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2871
timestamp 1666464484
transform 1 0 52976 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2872
timestamp 1666464484
transform 1 0 60928 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2873
timestamp 1666464484
transform 1 0 68880 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2874
timestamp 1666464484
transform 1 0 76832 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2875
timestamp 1666464484
transform 1 0 84784 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2876
timestamp 1666464484
transform 1 0 92736 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2877
timestamp 1666464484
transform 1 0 100688 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2878
timestamp 1666464484
transform 1 0 108640 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2879
timestamp 1666464484
transform 1 0 116592 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2880
timestamp 1666464484
transform 1 0 124544 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2881
timestamp 1666464484
transform 1 0 132496 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2882
timestamp 1666464484
transform 1 0 140448 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2883
timestamp 1666464484
transform 1 0 148400 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2884
timestamp 1666464484
transform 1 0 156352 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2885
timestamp 1666464484
transform 1 0 164304 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2886
timestamp 1666464484
transform 1 0 172256 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2887
timestamp 1666464484
transform 1 0 9296 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2888
timestamp 1666464484
transform 1 0 17248 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2889
timestamp 1666464484
transform 1 0 25200 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2890
timestamp 1666464484
transform 1 0 33152 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2891
timestamp 1666464484
transform 1 0 41104 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2892
timestamp 1666464484
transform 1 0 49056 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2893
timestamp 1666464484
transform 1 0 57008 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2894
timestamp 1666464484
transform 1 0 64960 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2895
timestamp 1666464484
transform 1 0 72912 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2896
timestamp 1666464484
transform 1 0 80864 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2897
timestamp 1666464484
transform 1 0 88816 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2898
timestamp 1666464484
transform 1 0 96768 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2899
timestamp 1666464484
transform 1 0 104720 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2900
timestamp 1666464484
transform 1 0 112672 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2901
timestamp 1666464484
transform 1 0 120624 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2902
timestamp 1666464484
transform 1 0 128576 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2903
timestamp 1666464484
transform 1 0 136528 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2904
timestamp 1666464484
transform 1 0 144480 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2905
timestamp 1666464484
transform 1 0 152432 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2906
timestamp 1666464484
transform 1 0 160384 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2907
timestamp 1666464484
transform 1 0 168336 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2908
timestamp 1666464484
transform 1 0 176288 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2909
timestamp 1666464484
transform 1 0 5264 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2910
timestamp 1666464484
transform 1 0 13216 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2911
timestamp 1666464484
transform 1 0 21168 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2912
timestamp 1666464484
transform 1 0 29120 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2913
timestamp 1666464484
transform 1 0 37072 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2914
timestamp 1666464484
transform 1 0 45024 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2915
timestamp 1666464484
transform 1 0 52976 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2916
timestamp 1666464484
transform 1 0 60928 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2917
timestamp 1666464484
transform 1 0 68880 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2918
timestamp 1666464484
transform 1 0 76832 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2919
timestamp 1666464484
transform 1 0 84784 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2920
timestamp 1666464484
transform 1 0 92736 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2921
timestamp 1666464484
transform 1 0 100688 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2922
timestamp 1666464484
transform 1 0 108640 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2923
timestamp 1666464484
transform 1 0 116592 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2924
timestamp 1666464484
transform 1 0 124544 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2925
timestamp 1666464484
transform 1 0 132496 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2926
timestamp 1666464484
transform 1 0 140448 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2927
timestamp 1666464484
transform 1 0 148400 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2928
timestamp 1666464484
transform 1 0 156352 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2929
timestamp 1666464484
transform 1 0 164304 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2930
timestamp 1666464484
transform 1 0 172256 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2931
timestamp 1666464484
transform 1 0 9296 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2932
timestamp 1666464484
transform 1 0 17248 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2933
timestamp 1666464484
transform 1 0 25200 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2934
timestamp 1666464484
transform 1 0 33152 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2935
timestamp 1666464484
transform 1 0 41104 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2936
timestamp 1666464484
transform 1 0 49056 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2937
timestamp 1666464484
transform 1 0 57008 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2938
timestamp 1666464484
transform 1 0 64960 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2939
timestamp 1666464484
transform 1 0 72912 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2940
timestamp 1666464484
transform 1 0 80864 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2941
timestamp 1666464484
transform 1 0 88816 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2942
timestamp 1666464484
transform 1 0 96768 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2943
timestamp 1666464484
transform 1 0 104720 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2944
timestamp 1666464484
transform 1 0 112672 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2945
timestamp 1666464484
transform 1 0 120624 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2946
timestamp 1666464484
transform 1 0 128576 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2947
timestamp 1666464484
transform 1 0 136528 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2948
timestamp 1666464484
transform 1 0 144480 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2949
timestamp 1666464484
transform 1 0 152432 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2950
timestamp 1666464484
transform 1 0 160384 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2951
timestamp 1666464484
transform 1 0 168336 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2952
timestamp 1666464484
transform 1 0 176288 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2953
timestamp 1666464484
transform 1 0 5264 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2954
timestamp 1666464484
transform 1 0 13216 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2955
timestamp 1666464484
transform 1 0 21168 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2956
timestamp 1666464484
transform 1 0 29120 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2957
timestamp 1666464484
transform 1 0 37072 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2958
timestamp 1666464484
transform 1 0 45024 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2959
timestamp 1666464484
transform 1 0 52976 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2960
timestamp 1666464484
transform 1 0 60928 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2961
timestamp 1666464484
transform 1 0 68880 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2962
timestamp 1666464484
transform 1 0 76832 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2963
timestamp 1666464484
transform 1 0 84784 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2964
timestamp 1666464484
transform 1 0 92736 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2965
timestamp 1666464484
transform 1 0 100688 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2966
timestamp 1666464484
transform 1 0 108640 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2967
timestamp 1666464484
transform 1 0 116592 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2968
timestamp 1666464484
transform 1 0 124544 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2969
timestamp 1666464484
transform 1 0 132496 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2970
timestamp 1666464484
transform 1 0 140448 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2971
timestamp 1666464484
transform 1 0 148400 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2972
timestamp 1666464484
transform 1 0 156352 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2973
timestamp 1666464484
transform 1 0 164304 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2974
timestamp 1666464484
transform 1 0 172256 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2975
timestamp 1666464484
transform 1 0 9296 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2976
timestamp 1666464484
transform 1 0 17248 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2977
timestamp 1666464484
transform 1 0 25200 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2978
timestamp 1666464484
transform 1 0 33152 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2979
timestamp 1666464484
transform 1 0 41104 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2980
timestamp 1666464484
transform 1 0 49056 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2981
timestamp 1666464484
transform 1 0 57008 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2982
timestamp 1666464484
transform 1 0 64960 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2983
timestamp 1666464484
transform 1 0 72912 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2984
timestamp 1666464484
transform 1 0 80864 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2985
timestamp 1666464484
transform 1 0 88816 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2986
timestamp 1666464484
transform 1 0 96768 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2987
timestamp 1666464484
transform 1 0 104720 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2988
timestamp 1666464484
transform 1 0 112672 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2989
timestamp 1666464484
transform 1 0 120624 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2990
timestamp 1666464484
transform 1 0 128576 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2991
timestamp 1666464484
transform 1 0 136528 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2992
timestamp 1666464484
transform 1 0 144480 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2993
timestamp 1666464484
transform 1 0 152432 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2994
timestamp 1666464484
transform 1 0 160384 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2995
timestamp 1666464484
transform 1 0 168336 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2996
timestamp 1666464484
transform 1 0 176288 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2997
timestamp 1666464484
transform 1 0 5264 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2998
timestamp 1666464484
transform 1 0 13216 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2999
timestamp 1666464484
transform 1 0 21168 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3000
timestamp 1666464484
transform 1 0 29120 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3001
timestamp 1666464484
transform 1 0 37072 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3002
timestamp 1666464484
transform 1 0 45024 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3003
timestamp 1666464484
transform 1 0 52976 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3004
timestamp 1666464484
transform 1 0 60928 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3005
timestamp 1666464484
transform 1 0 68880 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3006
timestamp 1666464484
transform 1 0 76832 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3007
timestamp 1666464484
transform 1 0 84784 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3008
timestamp 1666464484
transform 1 0 92736 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3009
timestamp 1666464484
transform 1 0 100688 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3010
timestamp 1666464484
transform 1 0 108640 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3011
timestamp 1666464484
transform 1 0 116592 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3012
timestamp 1666464484
transform 1 0 124544 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3013
timestamp 1666464484
transform 1 0 132496 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3014
timestamp 1666464484
transform 1 0 140448 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3015
timestamp 1666464484
transform 1 0 148400 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3016
timestamp 1666464484
transform 1 0 156352 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3017
timestamp 1666464484
transform 1 0 164304 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3018
timestamp 1666464484
transform 1 0 172256 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3019
timestamp 1666464484
transform 1 0 9296 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3020
timestamp 1666464484
transform 1 0 17248 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3021
timestamp 1666464484
transform 1 0 25200 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3022
timestamp 1666464484
transform 1 0 33152 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3023
timestamp 1666464484
transform 1 0 41104 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3024
timestamp 1666464484
transform 1 0 49056 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3025
timestamp 1666464484
transform 1 0 57008 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3026
timestamp 1666464484
transform 1 0 64960 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3027
timestamp 1666464484
transform 1 0 72912 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3028
timestamp 1666464484
transform 1 0 80864 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3029
timestamp 1666464484
transform 1 0 88816 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3030
timestamp 1666464484
transform 1 0 96768 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3031
timestamp 1666464484
transform 1 0 104720 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3032
timestamp 1666464484
transform 1 0 112672 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3033
timestamp 1666464484
transform 1 0 120624 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3034
timestamp 1666464484
transform 1 0 128576 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3035
timestamp 1666464484
transform 1 0 136528 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3036
timestamp 1666464484
transform 1 0 144480 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3037
timestamp 1666464484
transform 1 0 152432 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3038
timestamp 1666464484
transform 1 0 160384 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3039
timestamp 1666464484
transform 1 0 168336 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3040
timestamp 1666464484
transform 1 0 176288 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3041
timestamp 1666464484
transform 1 0 5264 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3042
timestamp 1666464484
transform 1 0 13216 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3043
timestamp 1666464484
transform 1 0 21168 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3044
timestamp 1666464484
transform 1 0 29120 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3045
timestamp 1666464484
transform 1 0 37072 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3046
timestamp 1666464484
transform 1 0 45024 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3047
timestamp 1666464484
transform 1 0 52976 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3048
timestamp 1666464484
transform 1 0 60928 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3049
timestamp 1666464484
transform 1 0 68880 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3050
timestamp 1666464484
transform 1 0 76832 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3051
timestamp 1666464484
transform 1 0 84784 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3052
timestamp 1666464484
transform 1 0 92736 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3053
timestamp 1666464484
transform 1 0 100688 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3054
timestamp 1666464484
transform 1 0 108640 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3055
timestamp 1666464484
transform 1 0 116592 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3056
timestamp 1666464484
transform 1 0 124544 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3057
timestamp 1666464484
transform 1 0 132496 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3058
timestamp 1666464484
transform 1 0 140448 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3059
timestamp 1666464484
transform 1 0 148400 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3060
timestamp 1666464484
transform 1 0 156352 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3061
timestamp 1666464484
transform 1 0 164304 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3062
timestamp 1666464484
transform 1 0 172256 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3063
timestamp 1666464484
transform 1 0 9296 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3064
timestamp 1666464484
transform 1 0 17248 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3065
timestamp 1666464484
transform 1 0 25200 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3066
timestamp 1666464484
transform 1 0 33152 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3067
timestamp 1666464484
transform 1 0 41104 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3068
timestamp 1666464484
transform 1 0 49056 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3069
timestamp 1666464484
transform 1 0 57008 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3070
timestamp 1666464484
transform 1 0 64960 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3071
timestamp 1666464484
transform 1 0 72912 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3072
timestamp 1666464484
transform 1 0 80864 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3073
timestamp 1666464484
transform 1 0 88816 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3074
timestamp 1666464484
transform 1 0 96768 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3075
timestamp 1666464484
transform 1 0 104720 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3076
timestamp 1666464484
transform 1 0 112672 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3077
timestamp 1666464484
transform 1 0 120624 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3078
timestamp 1666464484
transform 1 0 128576 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3079
timestamp 1666464484
transform 1 0 136528 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3080
timestamp 1666464484
transform 1 0 144480 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3081
timestamp 1666464484
transform 1 0 152432 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3082
timestamp 1666464484
transform 1 0 160384 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3083
timestamp 1666464484
transform 1 0 168336 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3084
timestamp 1666464484
transform 1 0 176288 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3085
timestamp 1666464484
transform 1 0 5264 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3086
timestamp 1666464484
transform 1 0 13216 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3087
timestamp 1666464484
transform 1 0 21168 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3088
timestamp 1666464484
transform 1 0 29120 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3089
timestamp 1666464484
transform 1 0 37072 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3090
timestamp 1666464484
transform 1 0 45024 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3091
timestamp 1666464484
transform 1 0 52976 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3092
timestamp 1666464484
transform 1 0 60928 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3093
timestamp 1666464484
transform 1 0 68880 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3094
timestamp 1666464484
transform 1 0 76832 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3095
timestamp 1666464484
transform 1 0 84784 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3096
timestamp 1666464484
transform 1 0 92736 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3097
timestamp 1666464484
transform 1 0 100688 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3098
timestamp 1666464484
transform 1 0 108640 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3099
timestamp 1666464484
transform 1 0 116592 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3100
timestamp 1666464484
transform 1 0 124544 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3101
timestamp 1666464484
transform 1 0 132496 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3102
timestamp 1666464484
transform 1 0 140448 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3103
timestamp 1666464484
transform 1 0 148400 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3104
timestamp 1666464484
transform 1 0 156352 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3105
timestamp 1666464484
transform 1 0 164304 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3106
timestamp 1666464484
transform 1 0 172256 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3107
timestamp 1666464484
transform 1 0 9296 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3108
timestamp 1666464484
transform 1 0 17248 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3109
timestamp 1666464484
transform 1 0 25200 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3110
timestamp 1666464484
transform 1 0 33152 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3111
timestamp 1666464484
transform 1 0 41104 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3112
timestamp 1666464484
transform 1 0 49056 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3113
timestamp 1666464484
transform 1 0 57008 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3114
timestamp 1666464484
transform 1 0 64960 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3115
timestamp 1666464484
transform 1 0 72912 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3116
timestamp 1666464484
transform 1 0 80864 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3117
timestamp 1666464484
transform 1 0 88816 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3118
timestamp 1666464484
transform 1 0 96768 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3119
timestamp 1666464484
transform 1 0 104720 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3120
timestamp 1666464484
transform 1 0 112672 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3121
timestamp 1666464484
transform 1 0 120624 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3122
timestamp 1666464484
transform 1 0 128576 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3123
timestamp 1666464484
transform 1 0 136528 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3124
timestamp 1666464484
transform 1 0 144480 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3125
timestamp 1666464484
transform 1 0 152432 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3126
timestamp 1666464484
transform 1 0 160384 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3127
timestamp 1666464484
transform 1 0 168336 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3128
timestamp 1666464484
transform 1 0 176288 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3129
timestamp 1666464484
transform 1 0 5264 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3130
timestamp 1666464484
transform 1 0 13216 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3131
timestamp 1666464484
transform 1 0 21168 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3132
timestamp 1666464484
transform 1 0 29120 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3133
timestamp 1666464484
transform 1 0 37072 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3134
timestamp 1666464484
transform 1 0 45024 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3135
timestamp 1666464484
transform 1 0 52976 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3136
timestamp 1666464484
transform 1 0 60928 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3137
timestamp 1666464484
transform 1 0 68880 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3138
timestamp 1666464484
transform 1 0 76832 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3139
timestamp 1666464484
transform 1 0 84784 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3140
timestamp 1666464484
transform 1 0 92736 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3141
timestamp 1666464484
transform 1 0 100688 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3142
timestamp 1666464484
transform 1 0 108640 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3143
timestamp 1666464484
transform 1 0 116592 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3144
timestamp 1666464484
transform 1 0 124544 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3145
timestamp 1666464484
transform 1 0 132496 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3146
timestamp 1666464484
transform 1 0 140448 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3147
timestamp 1666464484
transform 1 0 148400 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3148
timestamp 1666464484
transform 1 0 156352 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3149
timestamp 1666464484
transform 1 0 164304 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3150
timestamp 1666464484
transform 1 0 172256 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3151
timestamp 1666464484
transform 1 0 9296 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3152
timestamp 1666464484
transform 1 0 17248 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3153
timestamp 1666464484
transform 1 0 25200 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3154
timestamp 1666464484
transform 1 0 33152 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3155
timestamp 1666464484
transform 1 0 41104 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3156
timestamp 1666464484
transform 1 0 49056 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3157
timestamp 1666464484
transform 1 0 57008 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3158
timestamp 1666464484
transform 1 0 64960 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3159
timestamp 1666464484
transform 1 0 72912 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3160
timestamp 1666464484
transform 1 0 80864 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3161
timestamp 1666464484
transform 1 0 88816 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3162
timestamp 1666464484
transform 1 0 96768 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3163
timestamp 1666464484
transform 1 0 104720 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3164
timestamp 1666464484
transform 1 0 112672 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3165
timestamp 1666464484
transform 1 0 120624 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3166
timestamp 1666464484
transform 1 0 128576 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3167
timestamp 1666464484
transform 1 0 136528 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3168
timestamp 1666464484
transform 1 0 144480 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3169
timestamp 1666464484
transform 1 0 152432 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3170
timestamp 1666464484
transform 1 0 160384 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3171
timestamp 1666464484
transform 1 0 168336 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3172
timestamp 1666464484
transform 1 0 176288 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3173
timestamp 1666464484
transform 1 0 5264 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3174
timestamp 1666464484
transform 1 0 13216 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3175
timestamp 1666464484
transform 1 0 21168 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3176
timestamp 1666464484
transform 1 0 29120 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3177
timestamp 1666464484
transform 1 0 37072 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3178
timestamp 1666464484
transform 1 0 45024 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3179
timestamp 1666464484
transform 1 0 52976 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3180
timestamp 1666464484
transform 1 0 60928 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3181
timestamp 1666464484
transform 1 0 68880 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3182
timestamp 1666464484
transform 1 0 76832 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3183
timestamp 1666464484
transform 1 0 84784 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3184
timestamp 1666464484
transform 1 0 92736 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3185
timestamp 1666464484
transform 1 0 100688 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3186
timestamp 1666464484
transform 1 0 108640 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3187
timestamp 1666464484
transform 1 0 116592 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3188
timestamp 1666464484
transform 1 0 124544 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3189
timestamp 1666464484
transform 1 0 132496 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3190
timestamp 1666464484
transform 1 0 140448 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3191
timestamp 1666464484
transform 1 0 148400 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3192
timestamp 1666464484
transform 1 0 156352 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3193
timestamp 1666464484
transform 1 0 164304 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3194
timestamp 1666464484
transform 1 0 172256 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3195
timestamp 1666464484
transform 1 0 9296 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3196
timestamp 1666464484
transform 1 0 17248 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3197
timestamp 1666464484
transform 1 0 25200 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3198
timestamp 1666464484
transform 1 0 33152 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3199
timestamp 1666464484
transform 1 0 41104 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3200
timestamp 1666464484
transform 1 0 49056 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3201
timestamp 1666464484
transform 1 0 57008 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3202
timestamp 1666464484
transform 1 0 64960 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3203
timestamp 1666464484
transform 1 0 72912 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3204
timestamp 1666464484
transform 1 0 80864 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3205
timestamp 1666464484
transform 1 0 88816 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3206
timestamp 1666464484
transform 1 0 96768 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3207
timestamp 1666464484
transform 1 0 104720 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3208
timestamp 1666464484
transform 1 0 112672 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3209
timestamp 1666464484
transform 1 0 120624 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3210
timestamp 1666464484
transform 1 0 128576 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3211
timestamp 1666464484
transform 1 0 136528 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3212
timestamp 1666464484
transform 1 0 144480 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3213
timestamp 1666464484
transform 1 0 152432 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3214
timestamp 1666464484
transform 1 0 160384 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3215
timestamp 1666464484
transform 1 0 168336 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3216
timestamp 1666464484
transform 1 0 176288 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3217
timestamp 1666464484
transform 1 0 5264 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3218
timestamp 1666464484
transform 1 0 13216 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3219
timestamp 1666464484
transform 1 0 21168 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3220
timestamp 1666464484
transform 1 0 29120 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3221
timestamp 1666464484
transform 1 0 37072 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3222
timestamp 1666464484
transform 1 0 45024 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3223
timestamp 1666464484
transform 1 0 52976 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3224
timestamp 1666464484
transform 1 0 60928 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3225
timestamp 1666464484
transform 1 0 68880 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3226
timestamp 1666464484
transform 1 0 76832 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3227
timestamp 1666464484
transform 1 0 84784 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3228
timestamp 1666464484
transform 1 0 92736 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3229
timestamp 1666464484
transform 1 0 100688 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3230
timestamp 1666464484
transform 1 0 108640 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3231
timestamp 1666464484
transform 1 0 116592 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3232
timestamp 1666464484
transform 1 0 124544 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3233
timestamp 1666464484
transform 1 0 132496 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3234
timestamp 1666464484
transform 1 0 140448 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3235
timestamp 1666464484
transform 1 0 148400 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3236
timestamp 1666464484
transform 1 0 156352 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3237
timestamp 1666464484
transform 1 0 164304 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3238
timestamp 1666464484
transform 1 0 172256 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3239
timestamp 1666464484
transform 1 0 9296 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3240
timestamp 1666464484
transform 1 0 17248 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3241
timestamp 1666464484
transform 1 0 25200 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3242
timestamp 1666464484
transform 1 0 33152 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3243
timestamp 1666464484
transform 1 0 41104 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3244
timestamp 1666464484
transform 1 0 49056 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3245
timestamp 1666464484
transform 1 0 57008 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3246
timestamp 1666464484
transform 1 0 64960 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3247
timestamp 1666464484
transform 1 0 72912 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3248
timestamp 1666464484
transform 1 0 80864 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3249
timestamp 1666464484
transform 1 0 88816 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3250
timestamp 1666464484
transform 1 0 96768 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3251
timestamp 1666464484
transform 1 0 104720 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3252
timestamp 1666464484
transform 1 0 112672 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3253
timestamp 1666464484
transform 1 0 120624 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3254
timestamp 1666464484
transform 1 0 128576 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3255
timestamp 1666464484
transform 1 0 136528 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3256
timestamp 1666464484
transform 1 0 144480 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3257
timestamp 1666464484
transform 1 0 152432 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3258
timestamp 1666464484
transform 1 0 160384 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3259
timestamp 1666464484
transform 1 0 168336 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3260
timestamp 1666464484
transform 1 0 176288 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3261
timestamp 1666464484
transform 1 0 5264 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3262
timestamp 1666464484
transform 1 0 13216 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3263
timestamp 1666464484
transform 1 0 21168 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3264
timestamp 1666464484
transform 1 0 29120 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3265
timestamp 1666464484
transform 1 0 37072 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3266
timestamp 1666464484
transform 1 0 45024 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3267
timestamp 1666464484
transform 1 0 52976 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3268
timestamp 1666464484
transform 1 0 60928 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3269
timestamp 1666464484
transform 1 0 68880 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3270
timestamp 1666464484
transform 1 0 76832 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3271
timestamp 1666464484
transform 1 0 84784 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3272
timestamp 1666464484
transform 1 0 92736 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3273
timestamp 1666464484
transform 1 0 100688 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3274
timestamp 1666464484
transform 1 0 108640 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3275
timestamp 1666464484
transform 1 0 116592 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3276
timestamp 1666464484
transform 1 0 124544 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3277
timestamp 1666464484
transform 1 0 132496 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3278
timestamp 1666464484
transform 1 0 140448 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3279
timestamp 1666464484
transform 1 0 148400 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3280
timestamp 1666464484
transform 1 0 156352 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3281
timestamp 1666464484
transform 1 0 164304 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3282
timestamp 1666464484
transform 1 0 172256 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3283
timestamp 1666464484
transform 1 0 9296 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3284
timestamp 1666464484
transform 1 0 17248 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3285
timestamp 1666464484
transform 1 0 25200 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3286
timestamp 1666464484
transform 1 0 33152 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3287
timestamp 1666464484
transform 1 0 41104 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3288
timestamp 1666464484
transform 1 0 49056 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3289
timestamp 1666464484
transform 1 0 57008 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3290
timestamp 1666464484
transform 1 0 64960 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3291
timestamp 1666464484
transform 1 0 72912 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3292
timestamp 1666464484
transform 1 0 80864 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3293
timestamp 1666464484
transform 1 0 88816 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3294
timestamp 1666464484
transform 1 0 96768 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3295
timestamp 1666464484
transform 1 0 104720 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3296
timestamp 1666464484
transform 1 0 112672 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3297
timestamp 1666464484
transform 1 0 120624 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3298
timestamp 1666464484
transform 1 0 128576 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3299
timestamp 1666464484
transform 1 0 136528 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3300
timestamp 1666464484
transform 1 0 144480 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3301
timestamp 1666464484
transform 1 0 152432 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3302
timestamp 1666464484
transform 1 0 160384 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3303
timestamp 1666464484
transform 1 0 168336 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3304
timestamp 1666464484
transform 1 0 176288 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3305
timestamp 1666464484
transform 1 0 5264 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3306
timestamp 1666464484
transform 1 0 13216 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3307
timestamp 1666464484
transform 1 0 21168 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3308
timestamp 1666464484
transform 1 0 29120 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3309
timestamp 1666464484
transform 1 0 37072 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3310
timestamp 1666464484
transform 1 0 45024 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3311
timestamp 1666464484
transform 1 0 52976 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3312
timestamp 1666464484
transform 1 0 60928 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3313
timestamp 1666464484
transform 1 0 68880 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3314
timestamp 1666464484
transform 1 0 76832 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3315
timestamp 1666464484
transform 1 0 84784 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3316
timestamp 1666464484
transform 1 0 92736 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3317
timestamp 1666464484
transform 1 0 100688 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3318
timestamp 1666464484
transform 1 0 108640 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3319
timestamp 1666464484
transform 1 0 116592 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3320
timestamp 1666464484
transform 1 0 124544 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3321
timestamp 1666464484
transform 1 0 132496 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3322
timestamp 1666464484
transform 1 0 140448 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3323
timestamp 1666464484
transform 1 0 148400 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3324
timestamp 1666464484
transform 1 0 156352 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3325
timestamp 1666464484
transform 1 0 164304 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3326
timestamp 1666464484
transform 1 0 172256 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3327
timestamp 1666464484
transform 1 0 9296 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3328
timestamp 1666464484
transform 1 0 17248 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3329
timestamp 1666464484
transform 1 0 25200 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3330
timestamp 1666464484
transform 1 0 33152 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3331
timestamp 1666464484
transform 1 0 41104 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3332
timestamp 1666464484
transform 1 0 49056 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3333
timestamp 1666464484
transform 1 0 57008 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3334
timestamp 1666464484
transform 1 0 64960 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3335
timestamp 1666464484
transform 1 0 72912 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3336
timestamp 1666464484
transform 1 0 80864 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3337
timestamp 1666464484
transform 1 0 88816 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3338
timestamp 1666464484
transform 1 0 96768 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3339
timestamp 1666464484
transform 1 0 104720 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3340
timestamp 1666464484
transform 1 0 112672 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3341
timestamp 1666464484
transform 1 0 120624 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3342
timestamp 1666464484
transform 1 0 128576 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3343
timestamp 1666464484
transform 1 0 136528 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3344
timestamp 1666464484
transform 1 0 144480 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3345
timestamp 1666464484
transform 1 0 152432 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3346
timestamp 1666464484
transform 1 0 160384 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3347
timestamp 1666464484
transform 1 0 168336 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3348
timestamp 1666464484
transform 1 0 176288 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3349
timestamp 1666464484
transform 1 0 5264 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3350
timestamp 1666464484
transform 1 0 13216 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3351
timestamp 1666464484
transform 1 0 21168 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3352
timestamp 1666464484
transform 1 0 29120 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3353
timestamp 1666464484
transform 1 0 37072 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3354
timestamp 1666464484
transform 1 0 45024 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3355
timestamp 1666464484
transform 1 0 52976 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3356
timestamp 1666464484
transform 1 0 60928 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3357
timestamp 1666464484
transform 1 0 68880 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3358
timestamp 1666464484
transform 1 0 76832 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3359
timestamp 1666464484
transform 1 0 84784 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3360
timestamp 1666464484
transform 1 0 92736 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3361
timestamp 1666464484
transform 1 0 100688 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3362
timestamp 1666464484
transform 1 0 108640 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3363
timestamp 1666464484
transform 1 0 116592 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3364
timestamp 1666464484
transform 1 0 124544 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3365
timestamp 1666464484
transform 1 0 132496 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3366
timestamp 1666464484
transform 1 0 140448 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3367
timestamp 1666464484
transform 1 0 148400 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3368
timestamp 1666464484
transform 1 0 156352 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3369
timestamp 1666464484
transform 1 0 164304 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3370
timestamp 1666464484
transform 1 0 172256 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3371
timestamp 1666464484
transform 1 0 9296 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3372
timestamp 1666464484
transform 1 0 17248 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3373
timestamp 1666464484
transform 1 0 25200 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3374
timestamp 1666464484
transform 1 0 33152 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3375
timestamp 1666464484
transform 1 0 41104 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3376
timestamp 1666464484
transform 1 0 49056 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3377
timestamp 1666464484
transform 1 0 57008 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3378
timestamp 1666464484
transform 1 0 64960 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3379
timestamp 1666464484
transform 1 0 72912 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3380
timestamp 1666464484
transform 1 0 80864 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3381
timestamp 1666464484
transform 1 0 88816 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3382
timestamp 1666464484
transform 1 0 96768 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3383
timestamp 1666464484
transform 1 0 104720 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3384
timestamp 1666464484
transform 1 0 112672 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3385
timestamp 1666464484
transform 1 0 120624 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3386
timestamp 1666464484
transform 1 0 128576 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3387
timestamp 1666464484
transform 1 0 136528 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3388
timestamp 1666464484
transform 1 0 144480 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3389
timestamp 1666464484
transform 1 0 152432 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3390
timestamp 1666464484
transform 1 0 160384 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3391
timestamp 1666464484
transform 1 0 168336 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3392
timestamp 1666464484
transform 1 0 176288 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3393
timestamp 1666464484
transform 1 0 5264 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3394
timestamp 1666464484
transform 1 0 13216 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3395
timestamp 1666464484
transform 1 0 21168 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3396
timestamp 1666464484
transform 1 0 29120 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3397
timestamp 1666464484
transform 1 0 37072 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3398
timestamp 1666464484
transform 1 0 45024 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3399
timestamp 1666464484
transform 1 0 52976 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3400
timestamp 1666464484
transform 1 0 60928 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3401
timestamp 1666464484
transform 1 0 68880 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3402
timestamp 1666464484
transform 1 0 76832 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3403
timestamp 1666464484
transform 1 0 84784 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3404
timestamp 1666464484
transform 1 0 92736 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3405
timestamp 1666464484
transform 1 0 100688 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3406
timestamp 1666464484
transform 1 0 108640 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3407
timestamp 1666464484
transform 1 0 116592 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3408
timestamp 1666464484
transform 1 0 124544 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3409
timestamp 1666464484
transform 1 0 132496 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3410
timestamp 1666464484
transform 1 0 140448 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3411
timestamp 1666464484
transform 1 0 148400 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3412
timestamp 1666464484
transform 1 0 156352 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3413
timestamp 1666464484
transform 1 0 164304 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3414
timestamp 1666464484
transform 1 0 172256 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3415
timestamp 1666464484
transform 1 0 9296 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3416
timestamp 1666464484
transform 1 0 17248 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3417
timestamp 1666464484
transform 1 0 25200 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3418
timestamp 1666464484
transform 1 0 33152 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3419
timestamp 1666464484
transform 1 0 41104 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3420
timestamp 1666464484
transform 1 0 49056 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3421
timestamp 1666464484
transform 1 0 57008 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3422
timestamp 1666464484
transform 1 0 64960 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3423
timestamp 1666464484
transform 1 0 72912 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3424
timestamp 1666464484
transform 1 0 80864 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3425
timestamp 1666464484
transform 1 0 88816 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3426
timestamp 1666464484
transform 1 0 96768 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3427
timestamp 1666464484
transform 1 0 104720 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3428
timestamp 1666464484
transform 1 0 112672 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3429
timestamp 1666464484
transform 1 0 120624 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3430
timestamp 1666464484
transform 1 0 128576 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3431
timestamp 1666464484
transform 1 0 136528 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3432
timestamp 1666464484
transform 1 0 144480 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3433
timestamp 1666464484
transform 1 0 152432 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3434
timestamp 1666464484
transform 1 0 160384 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3435
timestamp 1666464484
transform 1 0 168336 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3436
timestamp 1666464484
transform 1 0 176288 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3437
timestamp 1666464484
transform 1 0 5264 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3438
timestamp 1666464484
transform 1 0 13216 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3439
timestamp 1666464484
transform 1 0 21168 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3440
timestamp 1666464484
transform 1 0 29120 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3441
timestamp 1666464484
transform 1 0 37072 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3442
timestamp 1666464484
transform 1 0 45024 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3443
timestamp 1666464484
transform 1 0 52976 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3444
timestamp 1666464484
transform 1 0 60928 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3445
timestamp 1666464484
transform 1 0 68880 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3446
timestamp 1666464484
transform 1 0 76832 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3447
timestamp 1666464484
transform 1 0 84784 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3448
timestamp 1666464484
transform 1 0 92736 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3449
timestamp 1666464484
transform 1 0 100688 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3450
timestamp 1666464484
transform 1 0 108640 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3451
timestamp 1666464484
transform 1 0 116592 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3452
timestamp 1666464484
transform 1 0 124544 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3453
timestamp 1666464484
transform 1 0 132496 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3454
timestamp 1666464484
transform 1 0 140448 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3455
timestamp 1666464484
transform 1 0 148400 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3456
timestamp 1666464484
transform 1 0 156352 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3457
timestamp 1666464484
transform 1 0 164304 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3458
timestamp 1666464484
transform 1 0 172256 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3459
timestamp 1666464484
transform 1 0 9296 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3460
timestamp 1666464484
transform 1 0 17248 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3461
timestamp 1666464484
transform 1 0 25200 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3462
timestamp 1666464484
transform 1 0 33152 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3463
timestamp 1666464484
transform 1 0 41104 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3464
timestamp 1666464484
transform 1 0 49056 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3465
timestamp 1666464484
transform 1 0 57008 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3466
timestamp 1666464484
transform 1 0 64960 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3467
timestamp 1666464484
transform 1 0 72912 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3468
timestamp 1666464484
transform 1 0 80864 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3469
timestamp 1666464484
transform 1 0 88816 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3470
timestamp 1666464484
transform 1 0 96768 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3471
timestamp 1666464484
transform 1 0 104720 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3472
timestamp 1666464484
transform 1 0 112672 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3473
timestamp 1666464484
transform 1 0 120624 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3474
timestamp 1666464484
transform 1 0 128576 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3475
timestamp 1666464484
transform 1 0 136528 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3476
timestamp 1666464484
transform 1 0 144480 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3477
timestamp 1666464484
transform 1 0 152432 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3478
timestamp 1666464484
transform 1 0 160384 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3479
timestamp 1666464484
transform 1 0 168336 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3480
timestamp 1666464484
transform 1 0 176288 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3481
timestamp 1666464484
transform 1 0 5264 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3482
timestamp 1666464484
transform 1 0 9184 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3483
timestamp 1666464484
transform 1 0 13104 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3484
timestamp 1666464484
transform 1 0 17024 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3485
timestamp 1666464484
transform 1 0 20944 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3486
timestamp 1666464484
transform 1 0 24864 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3487
timestamp 1666464484
transform 1 0 28784 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3488
timestamp 1666464484
transform 1 0 32704 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3489
timestamp 1666464484
transform 1 0 36624 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3490
timestamp 1666464484
transform 1 0 40544 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3491
timestamp 1666464484
transform 1 0 44464 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3492
timestamp 1666464484
transform 1 0 48384 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3493
timestamp 1666464484
transform 1 0 52304 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3494
timestamp 1666464484
transform 1 0 56224 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3495
timestamp 1666464484
transform 1 0 60144 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3496
timestamp 1666464484
transform 1 0 64064 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3497
timestamp 1666464484
transform 1 0 67984 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3498
timestamp 1666464484
transform 1 0 71904 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3499
timestamp 1666464484
transform 1 0 75824 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3500
timestamp 1666464484
transform 1 0 79744 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3501
timestamp 1666464484
transform 1 0 83664 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3502
timestamp 1666464484
transform 1 0 87584 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3503
timestamp 1666464484
transform 1 0 91504 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3504
timestamp 1666464484
transform 1 0 95424 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3505
timestamp 1666464484
transform 1 0 99344 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3506
timestamp 1666464484
transform 1 0 103264 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3507
timestamp 1666464484
transform 1 0 107184 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3508
timestamp 1666464484
transform 1 0 111104 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3509
timestamp 1666464484
transform 1 0 115024 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3510
timestamp 1666464484
transform 1 0 118944 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3511
timestamp 1666464484
transform 1 0 122864 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3512
timestamp 1666464484
transform 1 0 126784 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3513
timestamp 1666464484
transform 1 0 130704 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3514
timestamp 1666464484
transform 1 0 134624 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3515
timestamp 1666464484
transform 1 0 138544 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3516
timestamp 1666464484
transform 1 0 142464 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3517
timestamp 1666464484
transform 1 0 146384 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3518
timestamp 1666464484
transform 1 0 150304 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3519
timestamp 1666464484
transform 1 0 154224 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3520
timestamp 1666464484
transform 1 0 158144 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3521
timestamp 1666464484
transform 1 0 162064 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3522
timestamp 1666464484
transform 1 0 165984 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3523
timestamp 1666464484
transform 1 0 169904 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3524
timestamp 1666464484
transform 1 0 173824 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_3525
timestamp 1666464484
transform 1 0 177744 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _346_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 89152 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _347_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 8288 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _348_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 135856 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _349_
timestamp 1666464484
transform -1 0 134848 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _350_
timestamp 1666464484
transform 1 0 132496 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _351_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 92848 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _352_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 64624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _353_
timestamp 1666464484
transform 1 0 55216 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _354_
timestamp 1666464484
transform -1 0 42000 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _355_
timestamp 1666464484
transform -1 0 39200 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _356_
timestamp 1666464484
transform 1 0 103488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _357_
timestamp 1666464484
transform -1 0 116256 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _358_
timestamp 1666464484
transform -1 0 121632 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _359_
timestamp 1666464484
transform 1 0 128800 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _360_
timestamp 1666464484
transform -1 0 129584 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _361_
timestamp 1666464484
transform 1 0 128912 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _362_
timestamp 1666464484
transform -1 0 126000 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _363_
timestamp 1666464484
transform 1 0 123648 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _364_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 123312 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _365_
timestamp 1666464484
transform 1 0 140784 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _366_
timestamp 1666464484
transform -1 0 145488 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _367_
timestamp 1666464484
transform 1 0 92624 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _368_
timestamp 1666464484
transform 1 0 121856 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _369_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 113008 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _370_
timestamp 1666464484
transform 1 0 131488 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _371_
timestamp 1666464484
transform 1 0 138992 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _372_
timestamp 1666464484
transform 1 0 131600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _373_
timestamp 1666464484
transform 1 0 130704 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _374_
timestamp 1666464484
transform -1 0 128464 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _375_
timestamp 1666464484
transform 1 0 129808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _376_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 130368 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _377_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 128576 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _378_
timestamp 1666464484
transform -1 0 126224 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _379_
timestamp 1666464484
transform 1 0 140560 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _380_
timestamp 1666464484
transform 1 0 135632 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _381_
timestamp 1666464484
transform 1 0 146608 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _382_
timestamp 1666464484
transform -1 0 140000 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _383_
timestamp 1666464484
transform 1 0 139664 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _384_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 136416 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _385_
timestamp 1666464484
transform 1 0 147504 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _386_
timestamp 1666464484
transform -1 0 146384 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _387_
timestamp 1666464484
transform 1 0 148512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _388_
timestamp 1666464484
transform 1 0 148624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _389_
timestamp 1666464484
transform -1 0 145824 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _390_
timestamp 1666464484
transform -1 0 134960 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _391_
timestamp 1666464484
transform 1 0 137984 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _392_
timestamp 1666464484
transform 1 0 147728 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _393_
timestamp 1666464484
transform -1 0 130480 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _394_
timestamp 1666464484
transform 1 0 146832 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _395_
timestamp 1666464484
transform -1 0 134064 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _396_
timestamp 1666464484
transform 1 0 132832 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _397_
timestamp 1666464484
transform 1 0 142800 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _398_
timestamp 1666464484
transform 1 0 143808 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _399_
timestamp 1666464484
transform 1 0 144816 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _400_
timestamp 1666464484
transform -1 0 136192 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _401_
timestamp 1666464484
transform 1 0 141456 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _402_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 138768 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _403_
timestamp 1666464484
transform -1 0 124320 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1666464484
transform -1 0 92624 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _405_
timestamp 1666464484
transform 1 0 13888 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _406_
timestamp 1666464484
transform 1 0 39200 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _407_
timestamp 1666464484
transform 1 0 74704 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _408_
timestamp 1666464484
transform 1 0 75152 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_
timestamp 1666464484
transform -1 0 75712 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _410_
timestamp 1666464484
transform 1 0 63952 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _411_
timestamp 1666464484
transform 1 0 65296 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _412_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 67088 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _413_
timestamp 1666464484
transform 1 0 39424 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _414_
timestamp 1666464484
transform 1 0 40320 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _415_
timestamp 1666464484
transform 1 0 39984 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _416_
timestamp 1666464484
transform -1 0 59808 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _417_
timestamp 1666464484
transform 1 0 73808 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _418_
timestamp 1666464484
transform -1 0 73920 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _419_
timestamp 1666464484
transform 1 0 62160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _420_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 65744 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _421_
timestamp 1666464484
transform 1 0 78288 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _422_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 42112 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _423_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 67312 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _424_
timestamp 1666464484
transform -1 0 67312 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _425_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 67536 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _426_
timestamp 1666464484
transform -1 0 79632 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _427_
timestamp 1666464484
transform -1 0 66864 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _428_
timestamp 1666464484
transform 1 0 77504 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _429_
timestamp 1666464484
transform 1 0 42224 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _430_
timestamp 1666464484
transform 1 0 69216 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _431_
timestamp 1666464484
transform -1 0 69104 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _432_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 67312 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _433_
timestamp 1666464484
transform 1 0 42224 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _434_
timestamp 1666464484
transform 1 0 68320 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _435_
timestamp 1666464484
transform -1 0 68208 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _436_
timestamp 1666464484
transform -1 0 131376 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _437_
timestamp 1666464484
transform -1 0 128240 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _438_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 23856 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _439_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 65856 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _440_
timestamp 1666464484
transform 1 0 69776 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _441_
timestamp 1666464484
transform 1 0 76048 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _442_
timestamp 1666464484
transform 1 0 76832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _443_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 71008 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _444_
timestamp 1666464484
transform -1 0 72016 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _445_
timestamp 1666464484
transform -1 0 78064 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _446_
timestamp 1666464484
transform 1 0 70560 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _447_
timestamp 1666464484
transform 1 0 71232 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _448_
timestamp 1666464484
transform 1 0 73248 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _449_
timestamp 1666464484
transform 1 0 75040 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _450_
timestamp 1666464484
transform 1 0 70672 0 1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _451_
timestamp 1666464484
transform 1 0 71344 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _452_
timestamp 1666464484
transform 1 0 73248 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _453_
timestamp 1666464484
transform -1 0 74144 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _454_
timestamp 1666464484
transform 1 0 135296 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _455_
timestamp 1666464484
transform -1 0 134176 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _456_
timestamp 1666464484
transform 1 0 78624 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _457_
timestamp 1666464484
transform -1 0 76720 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _458_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 71792 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _459_
timestamp 1666464484
transform 1 0 75936 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _460_
timestamp 1666464484
transform 1 0 77168 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _461_
timestamp 1666464484
transform -1 0 76720 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _462_
timestamp 1666464484
transform 1 0 14784 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _463_
timestamp 1666464484
transform 1 0 80192 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _464_
timestamp 1666464484
transform 1 0 81984 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _465_
timestamp 1666464484
transform -1 0 87024 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _466_
timestamp 1666464484
transform 1 0 78064 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _467_
timestamp 1666464484
transform 1 0 80304 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _468_
timestamp 1666464484
transform 1 0 80752 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _469_
timestamp 1666464484
transform -1 0 84672 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _470_
timestamp 1666464484
transform 1 0 83104 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _471_
timestamp 1666464484
transform -1 0 78960 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _472_
timestamp 1666464484
transform 1 0 80640 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _473_
timestamp 1666464484
transform 1 0 75264 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _474_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 77168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _475_
timestamp 1666464484
transform -1 0 82656 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _476_
timestamp 1666464484
transform 1 0 84112 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _477_
timestamp 1666464484
transform 1 0 85120 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _478_
timestamp 1666464484
transform -1 0 102928 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _479_
timestamp 1666464484
transform -1 0 86016 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _480_
timestamp 1666464484
transform 1 0 82096 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _481_
timestamp 1666464484
transform 1 0 82096 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _482_
timestamp 1666464484
transform 1 0 84224 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _483_
timestamp 1666464484
transform -1 0 84112 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _484_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 51968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _485_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 76272 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _486_
timestamp 1666464484
transform 1 0 86128 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _487_
timestamp 1666464484
transform 1 0 85344 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _488_
timestamp 1666464484
transform 1 0 86240 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _489_
timestamp 1666464484
transform -1 0 86688 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _490_
timestamp 1666464484
transform 1 0 87136 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _491_
timestamp 1666464484
transform 1 0 89264 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _492_
timestamp 1666464484
transform 1 0 89600 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _493_
timestamp 1666464484
transform -1 0 87920 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _494_
timestamp 1666464484
transform 1 0 89152 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _495_
timestamp 1666464484
transform 1 0 89824 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _496_
timestamp 1666464484
transform 1 0 89824 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _497_
timestamp 1666464484
transform -1 0 88704 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _498_
timestamp 1666464484
transform 1 0 81648 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _499_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 68096 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _500_
timestamp 1666464484
transform -1 0 85792 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _501_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 82768 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _502_
timestamp 1666464484
transform -1 0 82992 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _503_
timestamp 1666464484
transform -1 0 144368 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _504_
timestamp 1666464484
transform 1 0 142688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _505_
timestamp 1666464484
transform 1 0 82768 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _506_
timestamp 1666464484
transform -1 0 83888 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _507_
timestamp 1666464484
transform -1 0 76720 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _508_
timestamp 1666464484
transform 1 0 88592 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _509_
timestamp 1666464484
transform 1 0 90160 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _510_
timestamp 1666464484
transform -1 0 91504 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _511_
timestamp 1666464484
transform 1 0 134400 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _512_
timestamp 1666464484
transform 1 0 16464 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _513_
timestamp 1666464484
transform -1 0 79520 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _514_
timestamp 1666464484
transform 1 0 74368 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _515_
timestamp 1666464484
transform 1 0 116928 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _516_
timestamp 1666464484
transform -1 0 92064 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _517_
timestamp 1666464484
transform 1 0 105168 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _518_
timestamp 1666464484
transform 1 0 78288 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _519_
timestamp 1666464484
transform 1 0 115136 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _520_
timestamp 1666464484
transform 1 0 117152 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _521_
timestamp 1666464484
transform -1 0 104608 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _522_
timestamp 1666464484
transform 1 0 117488 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _523_
timestamp 1666464484
transform -1 0 107632 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _524_
timestamp 1666464484
transform 1 0 81424 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _525_
timestamp 1666464484
transform 1 0 83328 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _526_
timestamp 1666464484
transform 1 0 117152 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _527_
timestamp 1666464484
transform 1 0 118160 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _528_
timestamp 1666464484
transform 1 0 119280 0 -1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _529_
timestamp 1666464484
transform -1 0 105728 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _530_
timestamp 1666464484
transform 1 0 116144 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _531_
timestamp 1666464484
transform 1 0 111888 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _532_
timestamp 1666464484
transform 1 0 119168 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _533_
timestamp 1666464484
transform 1 0 115024 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _534_
timestamp 1666464484
transform 1 0 120512 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _535_
timestamp 1666464484
transform -1 0 119616 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _536_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 119280 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _537_
timestamp 1666464484
transform -1 0 118944 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _538_
timestamp 1666464484
transform -1 0 120176 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _539_
timestamp 1666464484
transform 1 0 119056 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _540_
timestamp 1666464484
transform -1 0 118944 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _541_
timestamp 1666464484
transform 1 0 119952 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _542_
timestamp 1666464484
transform 1 0 120960 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _543_
timestamp 1666464484
transform -1 0 118720 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _544_
timestamp 1666464484
transform -1 0 119504 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _545_
timestamp 1666464484
transform 1 0 103824 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _546_
timestamp 1666464484
transform 1 0 104944 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _547_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 116480 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _548_
timestamp 1666464484
transform 1 0 121072 0 1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _549_
timestamp 1666464484
transform -1 0 116144 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _550_
timestamp 1666464484
transform 1 0 110992 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _551_
timestamp 1666464484
transform 1 0 113456 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _552_
timestamp 1666464484
transform 1 0 115360 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _553_
timestamp 1666464484
transform 1 0 116928 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _554_
timestamp 1666464484
transform -1 0 108528 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _555_
timestamp 1666464484
transform 1 0 142240 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _556_
timestamp 1666464484
transform 1 0 110992 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _557_
timestamp 1666464484
transform 1 0 111888 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _558_
timestamp 1666464484
transform 1 0 113008 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _559_
timestamp 1666464484
transform -1 0 110768 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _560_
timestamp 1666464484
transform 1 0 18592 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _561_
timestamp 1666464484
transform 1 0 79520 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _562_
timestamp 1666464484
transform 1 0 81200 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _563_
timestamp 1666464484
transform 1 0 98784 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _564_
timestamp 1666464484
transform -1 0 108304 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _565_
timestamp 1666464484
transform 1 0 107072 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _566_
timestamp 1666464484
transform 1 0 79856 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _567_
timestamp 1666464484
transform 1 0 94528 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _568_
timestamp 1666464484
transform 1 0 108080 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _569_
timestamp 1666464484
transform 1 0 108976 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _570_
timestamp 1666464484
transform 1 0 129584 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _571_
timestamp 1666464484
transform -1 0 98672 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _572_
timestamp 1666464484
transform -1 0 101360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _573_
timestamp 1666464484
transform -1 0 106064 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _574_
timestamp 1666464484
transform -1 0 97664 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _575_
timestamp 1666464484
transform 1 0 104048 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _576_
timestamp 1666464484
transform 1 0 102816 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _577_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 102928 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _578_
timestamp 1666464484
transform -1 0 102928 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _579_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 102256 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _580_
timestamp 1666464484
transform 1 0 101472 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _581_
timestamp 1666464484
transform 1 0 103152 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _582_
timestamp 1666464484
transform 1 0 101360 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _583_
timestamp 1666464484
transform 1 0 101920 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _584_
timestamp 1666464484
transform 1 0 105168 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _585_
timestamp 1666464484
transform -1 0 105504 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _586_
timestamp 1666464484
transform -1 0 97104 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _587_
timestamp 1666464484
transform -1 0 97888 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _588_
timestamp 1666464484
transform 1 0 95536 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _589_
timestamp 1666464484
transform 1 0 95760 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _590_
timestamp 1666464484
transform -1 0 159376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _591_
timestamp 1666464484
transform -1 0 137760 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _592_
timestamp 1666464484
transform -1 0 96656 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _593_
timestamp 1666464484
transform -1 0 95984 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _594_
timestamp 1666464484
transform 1 0 129808 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _595_
timestamp 1666464484
transform -1 0 98560 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _596_
timestamp 1666464484
transform 1 0 96656 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _597_
timestamp 1666464484
transform -1 0 92176 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _598_
timestamp 1666464484
transform 1 0 97664 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _599_
timestamp 1666464484
transform 1 0 97776 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _600_
timestamp 1666464484
transform 1 0 98448 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _601_
timestamp 1666464484
transform -1 0 99568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _602_
timestamp 1666464484
transform 1 0 98784 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _603_
timestamp 1666464484
transform -1 0 97552 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _604_
timestamp 1666464484
transform -1 0 95872 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _605_
timestamp 1666464484
transform -1 0 97552 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _606_
timestamp 1666464484
transform 1 0 96096 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _607_
timestamp 1666464484
transform 1 0 99120 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _608_
timestamp 1666464484
transform 1 0 101584 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _609_
timestamp 1666464484
transform -1 0 102144 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _610_
timestamp 1666464484
transform -1 0 98560 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _611_
timestamp 1666464484
transform 1 0 94976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _612_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 94640 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _613_
timestamp 1666464484
transform 1 0 95872 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _614_
timestamp 1666464484
transform 1 0 130480 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _615_
timestamp 1666464484
transform 1 0 99680 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _616_
timestamp 1666464484
transform -1 0 100240 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _617_
timestamp 1666464484
transform -1 0 44912 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _618_
timestamp 1666464484
transform 1 0 35616 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _619_
timestamp 1666464484
transform -1 0 38304 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _620_
timestamp 1666464484
transform 1 0 62384 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _621_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 62944 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _622_
timestamp 1666464484
transform 1 0 59248 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _623_
timestamp 1666464484
transform -1 0 49168 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _624_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 23408 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _625_
timestamp 1666464484
transform 1 0 14000 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _626_
timestamp 1666464484
transform -1 0 13104 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _627_
timestamp 1666464484
transform 1 0 17584 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _628_
timestamp 1666464484
transform -1 0 17136 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _629_
timestamp 1666464484
transform 1 0 19376 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _630_
timestamp 1666464484
transform -1 0 19824 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _631_
timestamp 1666464484
transform 1 0 21280 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _632_
timestamp 1666464484
transform -1 0 20832 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _633_
timestamp 1666464484
transform -1 0 31248 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _634_
timestamp 1666464484
transform 1 0 26432 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _635_
timestamp 1666464484
transform 1 0 25648 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _636_
timestamp 1666464484
transform -1 0 39648 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _637_
timestamp 1666464484
transform 1 0 37408 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _638_
timestamp 1666464484
transform 1 0 26096 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _639_
timestamp 1666464484
transform 1 0 25536 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _640_
timestamp 1666464484
transform 1 0 27216 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _641_
timestamp 1666464484
transform -1 0 27328 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _642_
timestamp 1666464484
transform 1 0 34608 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _643_
timestamp 1666464484
transform -1 0 36512 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _644_
timestamp 1666464484
transform 1 0 30128 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _645_
timestamp 1666464484
transform -1 0 30464 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _646_
timestamp 1666464484
transform 1 0 33936 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _647_
timestamp 1666464484
transform 1 0 33488 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _648_
timestamp 1666464484
transform -1 0 32368 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _649_
timestamp 1666464484
transform -1 0 35728 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _650_
timestamp 1666464484
transform -1 0 32480 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _651_
timestamp 1666464484
transform 1 0 45360 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _652_
timestamp 1666464484
transform -1 0 44128 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _653_
timestamp 1666464484
transform -1 0 45360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _654_
timestamp 1666464484
transform -1 0 48272 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _655_
timestamp 1666464484
transform -1 0 52864 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _656_
timestamp 1666464484
transform 1 0 53312 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _657_
timestamp 1666464484
transform 1 0 37632 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _658_
timestamp 1666464484
transform 1 0 37520 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _659_
timestamp 1666464484
transform 1 0 39536 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _660_
timestamp 1666464484
transform -1 0 39760 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _661_
timestamp 1666464484
transform 1 0 47712 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _662_
timestamp 1666464484
transform 1 0 45360 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _663_
timestamp 1666464484
transform 1 0 42336 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _664_
timestamp 1666464484
transform 1 0 44352 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _665_
timestamp 1666464484
transform -1 0 44240 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _666_
timestamp 1666464484
transform -1 0 51072 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _667_
timestamp 1666464484
transform -1 0 50624 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _668_
timestamp 1666464484
transform 1 0 47264 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _669_
timestamp 1666464484
transform -1 0 48160 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _670_
timestamp 1666464484
transform 1 0 45808 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _671_
timestamp 1666464484
transform -1 0 48160 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _672_
timestamp 1666464484
transform -1 0 51968 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _673_
timestamp 1666464484
transform -1 0 52640 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _674_
timestamp 1666464484
transform 1 0 54656 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _675_
timestamp 1666464484
transform 1 0 54096 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _676_
timestamp 1666464484
transform -1 0 54208 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _677_
timestamp 1666464484
transform 1 0 45360 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _678_
timestamp 1666464484
transform 1 0 56224 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _679_
timestamp 1666464484
transform -1 0 58240 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _680_
timestamp 1666464484
transform -1 0 56896 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _681_
timestamp 1666464484
transform -1 0 56448 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _682_
timestamp 1666464484
transform 1 0 57680 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _683_
timestamp 1666464484
transform -1 0 58016 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _684_
timestamp 1666464484
transform 1 0 60032 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _685_
timestamp 1666464484
transform 1 0 60032 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _686_
timestamp 1666464484
transform -1 0 60816 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _687_
timestamp 1666464484
transform -1 0 62048 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _688_
timestamp 1666464484
transform 1 0 63952 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _689_
timestamp 1666464484
transform 1 0 62160 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _690_
timestamp 1666464484
transform 1 0 63280 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _691_
timestamp 1666464484
transform 1 0 63280 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _692_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 38976 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _693_
timestamp 1666464484
transform 1 0 57568 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _694_
timestamp 1666464484
transform -1 0 66864 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _695_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 68656 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _696_
timestamp 1666464484
transform -1 0 69104 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _697_
timestamp 1666464484
transform -1 0 72800 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _698_
timestamp 1666464484
transform -1 0 72800 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _699_
timestamp 1666464484
transform 1 0 72464 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _700_
timestamp 1666464484
transform 1 0 75152 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _701_
timestamp 1666464484
transform -1 0 80080 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _702_
timestamp 1666464484
transform -1 0 86688 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _703_
timestamp 1666464484
transform -1 0 82544 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _704_
timestamp 1666464484
transform -1 0 88592 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _705_
timestamp 1666464484
transform 1 0 88144 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _706_
timestamp 1666464484
transform -1 0 92624 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _707_
timestamp 1666464484
transform 1 0 82544 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _708_
timestamp 1666464484
transform -1 0 92624 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _709_
timestamp 1666464484
transform 1 0 103264 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _710_
timestamp 1666464484
transform 1 0 105056 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _711_
timestamp 1666464484
transform 1 0 108976 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _712_
timestamp 1666464484
transform 1 0 109088 0 1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _713_
timestamp 1666464484
transform 1 0 108976 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _714_
timestamp 1666464484
transform 1 0 108976 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _715_
timestamp 1666464484
transform 1 0 108528 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _716_
timestamp 1666464484
transform 1 0 108976 0 -1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _717_
timestamp 1666464484
transform 1 0 109088 0 1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _718_
timestamp 1666464484
transform -1 0 104608 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _719_
timestamp 1666464484
transform 1 0 105056 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _720_
timestamp 1666464484
transform 1 0 94192 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _721_
timestamp 1666464484
transform -1 0 93408 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _722_
timestamp 1666464484
transform 1 0 98560 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _723_
timestamp 1666464484
transform 1 0 101024 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _724_
timestamp 1666464484
transform -1 0 100352 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _725_
timestamp 1666464484
transform -1 0 36176 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _726_
timestamp 1666464484
transform -1 0 61488 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _727_
timestamp 1666464484
transform 1 0 11872 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _728_
timestamp 1666464484
transform 1 0 15904 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _729_
timestamp 1666464484
transform 1 0 18032 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _730_
timestamp 1666464484
transform 1 0 19152 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _731_
timestamp 1666464484
transform 1 0 25536 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _732_
timestamp 1666464484
transform -1 0 38752 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _733_
timestamp 1666464484
transform -1 0 27216 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _734_
timestamp 1666464484
transform 1 0 25536 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _735_
timestamp 1666464484
transform -1 0 35168 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _736_
timestamp 1666464484
transform 1 0 29008 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _737_
timestamp 1666464484
transform 1 0 30464 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _738_
timestamp 1666464484
transform 1 0 30576 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _739_
timestamp 1666464484
transform -1 0 43568 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _740_
timestamp 1666464484
transform -1 0 52192 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _741_
timestamp 1666464484
transform 1 0 37408 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _742_
timestamp 1666464484
transform 1 0 37744 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _743_
timestamp 1666464484
transform 1 0 43232 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _744_
timestamp 1666464484
transform 1 0 42448 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _745_
timestamp 1666464484
transform -1 0 51296 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _746_
timestamp 1666464484
transform 1 0 46480 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _747_
timestamp 1666464484
transform -1 0 48608 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _748_
timestamp 1666464484
transform -1 0 52864 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _749_
timestamp 1666464484
transform 1 0 52304 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _750_
timestamp 1666464484
transform 1 0 53648 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _751_
timestamp 1666464484
transform 1 0 53312 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _752_
timestamp 1666464484
transform 1 0 56000 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _753_
timestamp 1666464484
transform -1 0 62608 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _754_
timestamp 1666464484
transform 1 0 57680 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _755_
timestamp 1666464484
transform 1 0 60368 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _756_
timestamp 1666464484
transform 1 0 62048 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _799_
timestamp 1666464484
transform -1 0 4928 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _800_
timestamp 1666464484
transform 1 0 7056 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _801_
timestamp 1666464484
transform 1 0 11536 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _802_
timestamp 1666464484
transform 1 0 16464 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _803_
timestamp 1666464484
transform 1 0 21280 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _804_
timestamp 1666464484
transform 1 0 25984 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _805_
timestamp 1666464484
transform 1 0 30688 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _806_
timestamp 1666464484
transform 1 0 35056 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _807_
timestamp 1666464484
transform 1 0 40096 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _808_
timestamp 1666464484
transform 1 0 44800 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _809_
timestamp 1666464484
transform 1 0 49504 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _810_
timestamp 1666464484
transform 1 0 54208 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _811_
timestamp 1666464484
transform 1 0 58576 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _812_
timestamp 1666464484
transform 1 0 63616 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _813_
timestamp 1666464484
transform 1 0 68320 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _814_
timestamp 1666464484
transform 1 0 73248 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _815_
timestamp 1666464484
transform 1 0 77728 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _816_
timestamp 1666464484
transform 1 0 82096 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _817_
timestamp 1666464484
transform -1 0 87808 0 1 114464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _818_
timestamp 1666464484
transform 1 0 91840 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _819_
timestamp 1666464484
transform -1 0 97776 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _820_
timestamp 1666464484
transform 1 0 101248 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _821_
timestamp 1666464484
transform 1 0 105840 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _822_
timestamp 1666464484
transform 1 0 110656 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _823_
timestamp 1666464484
transform 1 0 115360 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _824_
timestamp 1666464484
transform -1 0 121632 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _825_
timestamp 1666464484
transform 1 0 124656 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _826_
timestamp 1666464484
transform 1 0 129360 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _827_
timestamp 1666464484
transform 1 0 134176 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _828_
timestamp 1666464484
transform 1 0 138880 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _829_
timestamp 1666464484
transform 1 0 143584 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _830_
timestamp 1666464484
transform 1 0 148288 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _831_
timestamp 1666464484
transform 1 0 152992 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _832_
timestamp 1666464484
transform 1 0 157696 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _833_
timestamp 1666464484
transform 1 0 162400 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _834_
timestamp 1666464484
transform 1 0 167104 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _835_
timestamp 1666464484
transform 1 0 170464 0 -1 116032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _836_
timestamp 1666464484
transform 1 0 63056 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _837_
timestamp 1666464484
transform 1 0 65072 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _838_
timestamp 1666464484
transform 1 0 64176 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _839_
timestamp 1666464484
transform 1 0 67200 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _840_
timestamp 1666464484
transform -1 0 75712 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _841_
timestamp 1666464484
transform -1 0 74816 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _842_
timestamp 1666464484
transform 1 0 75152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _843_
timestamp 1666464484
transform 1 0 77168 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _844_
timestamp 1666464484
transform 1 0 78624 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _845_
timestamp 1666464484
transform 1 0 79744 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _846_
timestamp 1666464484
transform 1 0 81648 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _847_
timestamp 1666464484
transform 1 0 81872 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _848_
timestamp 1666464484
transform 1 0 86240 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _849_
timestamp 1666464484
transform -1 0 88928 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _850_
timestamp 1666464484
transform 1 0 87696 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _851_
timestamp 1666464484
transform 1 0 91616 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _852_
timestamp 1666464484
transform 1 0 93072 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _853_
timestamp 1666464484
transform 1 0 93968 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _854_
timestamp 1666464484
transform 1 0 94864 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _855_
timestamp 1666464484
transform -1 0 98784 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _856_
timestamp 1666464484
transform -1 0 100352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _857_
timestamp 1666464484
transform -1 0 103488 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _858_
timestamp 1666464484
transform -1 0 109648 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _859_
timestamp 1666464484
transform 1 0 103936 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _860_
timestamp 1666464484
transform 1 0 103936 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _861_
timestamp 1666464484
transform 1 0 107856 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _862_
timestamp 1666464484
transform 1 0 110096 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _863_
timestamp 1666464484
transform -1 0 113680 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _864_
timestamp 1666464484
transform 1 0 111888 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _865_
timestamp 1666464484
transform 1 0 114688 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _866_
timestamp 1666464484
transform 1 0 115248 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _867_
timestamp 1666464484
transform 1 0 117040 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 61264 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1666464484
transform -1 0 54992 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1666464484
transform -1 0 54992 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1666464484
transform 1 0 49392 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1666464484
transform 1 0 49392 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1666464484
transform 1 0 69216 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1666464484
transform 1 0 69216 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1666464484
transform 1 0 65296 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1666464484
transform 1 0 69216 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1666464484
transform -1 0 118832 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1666464484
transform -1 0 124768 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1666464484
transform -1 0 125104 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1666464484
transform -1 0 126896 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1666464484
transform -1 0 128688 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1666464484
transform -1 0 131712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1666464484
transform -1 0 133504 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1666464484
transform -1 0 134400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1666464484
transform -1 0 136528 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1666464484
transform -1 0 138320 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1666464484
transform -1 0 137536 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1666464484
transform -1 0 141344 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1666464484
transform -1 0 142240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1666464484
transform -1 0 142352 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1666464484
transform -1 0 145264 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1666464484
transform -1 0 146608 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1666464484
transform -1 0 148288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1666464484
transform -1 0 149408 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1666464484
transform -1 0 151312 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1666464484
transform -1 0 151760 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1666464484
transform -1 0 154000 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1666464484
transform -1 0 156128 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1666464484
transform -1 0 156800 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1666464484
transform -1 0 159152 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1666464484
transform -1 0 160944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1666464484
transform -1 0 161840 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1666464484
transform -1 0 163968 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1666464484
transform -1 0 165760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1666464484
transform -1 0 167888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1666464484
transform -1 0 169680 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1666464484
transform -1 0 170912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1666464484
transform -1 0 172704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1666464484
transform -1 0 123872 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1666464484
transform -1 0 125664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1666464484
transform -1 0 126560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1666464484
transform 1 0 127120 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1666464484
transform 1 0 128912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1666464484
transform 1 0 131936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1666464484
transform 1 0 132496 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1666464484
transform -1 0 135632 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1666464484
transform -1 0 137424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1666464484
transform 1 0 138880 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1666464484
transform -1 0 140448 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1666464484
transform -1 0 140896 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1666464484
transform -1 0 143472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1666464484
transform -1 0 144368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1666464484
transform -1 0 146160 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1666464484
transform -1 0 147392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1666464484
transform -1 0 150080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1666464484
transform -1 0 150192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1666464484
transform -1 0 152208 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1666464484
transform -1 0 153104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1666464484
transform -1 0 155232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1666464484
transform -1 0 157024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1666464484
transform -1 0 157920 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1666464484
transform -1 0 160048 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1666464484
transform -1 0 161840 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1666464484
transform -1 0 163072 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1666464484
transform -1 0 164864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1666464484
transform -1 0 166992 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1666464484
transform -1 0 168784 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1666464484
transform -1 0 169680 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1666464484
transform -1 0 171808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1666464484
transform -1 0 173600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  input65 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 6160 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1666464484
transform 1 0 7392 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1666464484
transform 1 0 9968 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input68
timestamp 1666464484
transform 1 0 29456 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input69
timestamp 1666464484
transform 1 0 28000 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input70
timestamp 1666464484
transform 1 0 29232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1666464484
transform 1 0 32368 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input72
timestamp 1666464484
transform 1 0 33712 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1666464484
transform 1 0 37408 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1666464484
transform 1 0 38640 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1666464484
transform 1 0 39536 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1666464484
transform 1 0 40432 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input77
timestamp 1666464484
transform 1 0 47152 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1666464484
transform 1 0 10976 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input79
timestamp 1666464484
transform 1 0 46256 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1666464484
transform 1 0 46368 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input81
timestamp 1666464484
transform 1 0 46816 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input82
timestamp 1666464484
transform 1 0 44240 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input83
timestamp 1666464484
transform 1 0 46368 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input84
timestamp 1666464484
transform 1 0 48720 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input85
timestamp 1666464484
transform 1 0 55216 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input86
timestamp 1666464484
transform 1 0 57568 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input87
timestamp 1666464484
transform 1 0 57344 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input88
timestamp 1666464484
transform 1 0 60256 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input89
timestamp 1666464484
transform 1 0 14448 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input90
timestamp 1666464484
transform 1 0 57344 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input91
timestamp 1666464484
transform 1 0 64848 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input92
timestamp 1666464484
transform 1 0 14112 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input93
timestamp 1666464484
transform 1 0 18256 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input94
timestamp 1666464484
transform 1 0 21056 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input95
timestamp 1666464484
transform 1 0 22288 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input96
timestamp 1666464484
transform 1 0 23968 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input97
timestamp 1666464484
transform 1 0 22624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input98
timestamp 1666464484
transform 1 0 25200 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input99
timestamp 1666464484
transform 1 0 11088 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input100
timestamp 1666464484
transform 1 0 12992 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input101
timestamp 1666464484
transform 1 0 15568 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input102
timestamp 1666464484
transform 1 0 15568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input103
timestamp 1666464484
transform -1 0 8960 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input104
timestamp 1666464484
transform 1 0 9408 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output105 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 4592 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output106
timestamp 1666464484
transform 1 0 50064 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output107
timestamp 1666464484
transform 1 0 54544 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output108
timestamp 1666464484
transform 1 0 59472 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output109
timestamp 1666464484
transform 1 0 64176 0 1 114464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output110
timestamp 1666464484
transform 1 0 68432 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output111
timestamp 1666464484
transform 1 0 73584 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output112
timestamp 1666464484
transform 1 0 78064 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output113
timestamp 1666464484
transform 1 0 82992 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output114
timestamp 1666464484
transform 1 0 87136 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output115
timestamp 1666464484
transform 1 0 92400 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output116
timestamp 1666464484
transform 1 0 7504 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output117
timestamp 1666464484
transform 1 0 97104 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output118
timestamp 1666464484
transform 1 0 101584 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output119
timestamp 1666464484
transform 1 0 107520 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output120
timestamp 1666464484
transform 1 0 111440 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output121
timestamp 1666464484
transform 1 0 115920 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output122
timestamp 1666464484
transform 1 0 120624 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output123
timestamp 1666464484
transform 1 0 125104 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output124
timestamp 1666464484
transform 1 0 131040 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output125
timestamp 1666464484
transform 1 0 134960 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output126
timestamp 1666464484
transform 1 0 139440 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output127
timestamp 1666464484
transform 1 0 12432 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output128
timestamp 1666464484
transform 1 0 144144 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output129
timestamp 1666464484
transform 1 0 148624 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output130
timestamp 1666464484
transform 1 0 154560 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output131
timestamp 1666464484
transform 1 0 158480 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output132
timestamp 1666464484
transform 1 0 162960 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output133
timestamp 1666464484
transform 1 0 167664 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output134
timestamp 1666464484
transform 1 0 172144 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output135
timestamp 1666464484
transform 1 0 17584 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output136
timestamp 1666464484
transform 1 0 21392 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output137
timestamp 1666464484
transform 1 0 26544 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output138
timestamp 1666464484
transform 1 0 31024 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output139
timestamp 1666464484
transform 1 0 35952 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output140
timestamp 1666464484
transform 1 0 41440 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output141
timestamp 1666464484
transform 1 0 44912 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output142
timestamp 1666464484
transform -1 0 7168 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output143
timestamp 1666464484
transform -1 0 54208 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output144
timestamp 1666464484
transform -1 0 58128 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output145
timestamp 1666464484
transform -1 0 62608 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output146
timestamp 1666464484
transform -1 0 67312 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output147
timestamp 1666464484
transform -1 0 71792 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output148
timestamp 1666464484
transform -1 0 77728 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output149
timestamp 1666464484
transform -1 0 81648 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output150
timestamp 1666464484
transform -1 0 86128 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output151
timestamp 1666464484
transform -1 0 90832 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output152
timestamp 1666464484
transform -1 0 95536 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output153
timestamp 1666464484
transform -1 0 11088 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output154
timestamp 1666464484
transform -1 0 101248 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output155
timestamp 1666464484
transform -1 0 105168 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output156
timestamp 1666464484
transform -1 0 109648 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output157
timestamp 1666464484
transform -1 0 114800 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output158
timestamp 1666464484
transform 1 0 117488 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output159
timestamp 1666464484
transform 1 0 123200 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output160
timestamp 1666464484
transform 1 0 127120 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output161
timestamp 1666464484
transform 1 0 131600 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output162
timestamp 1666464484
transform 1 0 136752 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output163
timestamp 1666464484
transform 1 0 141008 0 -1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output164
timestamp 1666464484
transform -1 0 15568 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output165
timestamp 1666464484
transform 1 0 146720 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output166
timestamp 1666464484
transform 1 0 150640 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output167
timestamp 1666464484
transform -1 0 20272 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output168
timestamp 1666464484
transform -1 0 24752 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output169
timestamp 1666464484
transform -1 0 30688 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output170
timestamp 1666464484
transform -1 0 34608 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output171
timestamp 1666464484
transform -1 0 39088 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output172
timestamp 1666464484
transform -1 0 43792 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output173
timestamp 1666464484
transform -1 0 48272 0 1 116032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output174
timestamp 1666464484
transform 1 0 65968 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output175
timestamp 1666464484
transform 1 0 81984 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output176
timestamp 1666464484
transform 1 0 84112 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output177
timestamp 1666464484
transform -1 0 87472 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output178
timestamp 1666464484
transform -1 0 88704 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output179
timestamp 1666464484
transform 1 0 89488 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output180
timestamp 1666464484
transform 1 0 91840 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output181
timestamp 1666464484
transform 1 0 93632 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output182
timestamp 1666464484
transform 1 0 94528 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output183
timestamp 1666464484
transform 1 0 96208 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output184
timestamp 1666464484
transform 1 0 97888 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output185
timestamp 1666464484
transform 1 0 68320 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output186
timestamp 1666464484
transform 1 0 99680 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output187
timestamp 1666464484
transform -1 0 103040 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output188
timestamp 1666464484
transform -1 0 105168 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output189
timestamp 1666464484
transform 1 0 105392 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output190
timestamp 1666464484
transform 1 0 106288 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output191
timestamp 1666464484
transform 1 0 107968 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output192
timestamp 1666464484
transform -1 0 111440 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output193
timestamp 1666464484
transform -1 0 113008 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output194
timestamp 1666464484
transform 1 0 113232 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output195
timestamp 1666464484
transform 1 0 115360 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output196
timestamp 1666464484
transform 1 0 69216 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output197
timestamp 1666464484
transform 1 0 117152 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output198
timestamp 1666464484
transform 1 0 119280 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output199
timestamp 1666464484
transform 1 0 70224 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output200
timestamp 1666464484
transform -1 0 73920 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output201
timestamp 1666464484
transform 1 0 74144 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output202
timestamp 1666464484
transform 1 0 76048 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output203
timestamp 1666464484
transform 1 0 77728 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output204
timestamp 1666464484
transform 1 0 79184 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output205
timestamp 1666464484
transform 1 0 80192 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output206
timestamp 1666464484
transform -1 0 8736 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output207
timestamp 1666464484
transform -1 0 11200 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output208
timestamp 1666464484
transform -1 0 31136 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output209
timestamp 1666464484
transform -1 0 32704 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output210
timestamp 1666464484
transform -1 0 34608 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output211
timestamp 1666464484
transform 1 0 33936 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output212
timestamp 1666464484
transform -1 0 36512 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output213
timestamp 1666464484
transform 1 0 37072 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output214
timestamp 1666464484
transform -1 0 40432 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output215
timestamp 1666464484
transform 1 0 40992 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output216
timestamp 1666464484
transform -1 0 44352 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output217
timestamp 1666464484
transform -1 0 45136 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output218
timestamp 1666464484
transform 1 0 11424 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output219
timestamp 1666464484
transform -1 0 46480 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output220
timestamp 1666464484
transform -1 0 48272 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output221
timestamp 1666464484
transform 1 0 46704 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output222
timestamp 1666464484
transform 1 0 51296 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output223
timestamp 1666464484
transform -1 0 54320 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output224
timestamp 1666464484
transform -1 0 56784 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output225
timestamp 1666464484
transform -1 0 56112 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output226
timestamp 1666464484
transform -1 0 58240 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output227
timestamp 1666464484
transform -1 0 60032 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output228
timestamp 1666464484
transform 1 0 60592 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output229
timestamp 1666464484
transform 1 0 15008 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output230
timestamp 1666464484
transform -1 0 63952 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output231
timestamp 1666464484
transform 1 0 65296 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output232
timestamp 1666464484
transform -1 0 18928 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output233
timestamp 1666464484
transform -1 0 21056 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output234
timestamp 1666464484
transform -1 0 20832 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output235
timestamp 1666464484
transform -1 0 23744 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output236
timestamp 1666464484
transform 1 0 23520 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output237
timestamp 1666464484
transform -1 0 24752 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output238
timestamp 1666464484
transform -1 0 29008 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_239 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 177520 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_240
timestamp 1666464484
transform -1 0 155568 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_241
timestamp 1666464484
transform -1 0 160720 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_242
timestamp 1666464484
transform -1 0 165200 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_243
timestamp 1666464484
transform -1 0 170688 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_244
timestamp 1666464484
transform -1 0 174608 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_245
timestamp 1666464484
transform 1 0 177856 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_246
timestamp 1666464484
transform -1 0 173376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_247
timestamp 1666464484
transform -1 0 174608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_248
timestamp 1666464484
transform -1 0 175280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_249
timestamp 1666464484
transform -1 0 122752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_250
timestamp 1666464484
transform -1 0 122752 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_251
timestamp 1666464484
transform -1 0 123424 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_252
timestamp 1666464484
transform -1 0 125216 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_253
timestamp 1666464484
transform -1 0 126896 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_254
timestamp 1666464484
transform -1 0 130144 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_255
timestamp 1666464484
transform -1 0 132048 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_256
timestamp 1666464484
transform -1 0 131936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_257
timestamp 1666464484
transform -1 0 133616 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_258
timestamp 1666464484
transform -1 0 135296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_259
timestamp 1666464484
transform -1 0 136976 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_260
timestamp 1666464484
transform -1 0 138656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_261
timestamp 1666464484
transform -1 0 140336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_262
timestamp 1666464484
transform -1 0 142016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_263
timestamp 1666464484
transform -1 0 143696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_264
timestamp 1666464484
transform -1 0 145376 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_265
timestamp 1666464484
transform -1 0 147056 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_266
timestamp 1666464484
transform -1 0 150864 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_267
timestamp 1666464484
transform -1 0 150416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_268
timestamp 1666464484
transform -1 0 152096 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_269
timestamp 1666464484
transform -1 0 153776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_270
timestamp 1666464484
transform -1 0 155456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_271
timestamp 1666464484
transform -1 0 157472 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_272
timestamp 1666464484
transform -1 0 158704 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_273
timestamp 1666464484
transform -1 0 160272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_274
timestamp 1666464484
transform -1 0 162512 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_275
timestamp 1666464484
transform -1 0 163856 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_276
timestamp 1666464484
transform -1 0 165536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_277
timestamp 1666464484
transform -1 0 167216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_278
timestamp 1666464484
transform 1 0 167776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_279
timestamp 1666464484
transform -1 0 170576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_280
timestamp 1666464484
transform -1 0 172256 0 -1 4704
box -86 -86 534 870
<< labels >>
flabel metal2 s 1344 119200 1456 120000 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 48384 119200 48496 120000 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 53088 119200 53200 120000 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 57792 119200 57904 120000 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 62496 119200 62608 120000 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 67200 119200 67312 120000 0 FreeSans 448 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 71904 119200 72016 120000 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 76608 119200 76720 120000 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 81312 119200 81424 120000 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 86016 119200 86128 120000 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 90720 119200 90832 120000 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 6048 119200 6160 120000 0 FreeSans 448 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 95424 119200 95536 120000 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 100128 119200 100240 120000 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 104832 119200 104944 120000 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 109536 119200 109648 120000 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 114240 119200 114352 120000 0 FreeSans 448 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 118944 119200 119056 120000 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 123648 119200 123760 120000 0 FreeSans 448 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 128352 119200 128464 120000 0 FreeSans 448 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 133056 119200 133168 120000 0 FreeSans 448 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 137760 119200 137872 120000 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 10752 119200 10864 120000 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 142464 119200 142576 120000 0 FreeSans 448 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 147168 119200 147280 120000 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 151872 119200 151984 120000 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 156576 119200 156688 120000 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 161280 119200 161392 120000 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 165984 119200 166096 120000 0 FreeSans 448 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 170688 119200 170800 120000 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 175392 119200 175504 120000 0 FreeSans 448 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 15456 119200 15568 120000 0 FreeSans 448 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 20160 119200 20272 120000 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 24864 119200 24976 120000 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 29568 119200 29680 120000 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 34272 119200 34384 120000 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 38976 119200 39088 120000 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 43680 119200 43792 120000 0 FreeSans 448 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 2912 119200 3024 120000 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 49952 119200 50064 120000 0 FreeSans 448 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 54656 119200 54768 120000 0 FreeSans 448 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 59360 119200 59472 120000 0 FreeSans 448 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 64064 119200 64176 120000 0 FreeSans 448 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 68768 119200 68880 120000 0 FreeSans 448 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 73472 119200 73584 120000 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 78176 119200 78288 120000 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 82880 119200 82992 120000 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 87584 119200 87696 120000 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 92288 119200 92400 120000 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 7616 119200 7728 120000 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 96992 119200 97104 120000 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 101696 119200 101808 120000 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 106400 119200 106512 120000 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 111104 119200 111216 120000 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 115808 119200 115920 120000 0 FreeSans 448 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 120512 119200 120624 120000 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 125216 119200 125328 120000 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 129920 119200 130032 120000 0 FreeSans 448 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 134624 119200 134736 120000 0 FreeSans 448 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 139328 119200 139440 120000 0 FreeSans 448 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 12320 119200 12432 120000 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 144032 119200 144144 120000 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 148736 119200 148848 120000 0 FreeSans 448 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 153440 119200 153552 120000 0 FreeSans 448 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 158144 119200 158256 120000 0 FreeSans 448 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 162848 119200 162960 120000 0 FreeSans 448 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 167552 119200 167664 120000 0 FreeSans 448 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 172256 119200 172368 120000 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 176960 119200 177072 120000 0 FreeSans 448 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 17024 119200 17136 120000 0 FreeSans 448 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 21728 119200 21840 120000 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 26432 119200 26544 120000 0 FreeSans 448 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 31136 119200 31248 120000 0 FreeSans 448 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 35840 119200 35952 120000 0 FreeSans 448 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 40544 119200 40656 120000 0 FreeSans 448 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 45248 119200 45360 120000 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 4480 119200 4592 120000 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 51520 119200 51632 120000 0 FreeSans 448 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 56224 119200 56336 120000 0 FreeSans 448 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 60928 119200 61040 120000 0 FreeSans 448 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 65632 119200 65744 120000 0 FreeSans 448 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 70336 119200 70448 120000 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 75040 119200 75152 120000 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 79744 119200 79856 120000 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 84448 119200 84560 120000 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 89152 119200 89264 120000 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 93856 119200 93968 120000 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 9184 119200 9296 120000 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 98560 119200 98672 120000 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 103264 119200 103376 120000 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 107968 119200 108080 120000 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 112672 119200 112784 120000 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 117376 119200 117488 120000 0 FreeSans 448 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 122080 119200 122192 120000 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 126784 119200 126896 120000 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 131488 119200 131600 120000 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 136192 119200 136304 120000 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 140896 119200 141008 120000 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 13888 119200 14000 120000 0 FreeSans 448 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 145600 119200 145712 120000 0 FreeSans 448 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 150304 119200 150416 120000 0 FreeSans 448 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 155008 119200 155120 120000 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 159712 119200 159824 120000 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 164416 119200 164528 120000 0 FreeSans 448 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 169120 119200 169232 120000 0 FreeSans 448 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 173824 119200 173936 120000 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 178528 119200 178640 120000 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 18592 119200 18704 120000 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 23296 119200 23408 120000 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 28000 119200 28112 120000 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 32704 119200 32816 120000 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 37408 119200 37520 120000 0 FreeSans 448 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 42112 119200 42224 120000 0 FreeSans 448 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 46816 119200 46928 120000 0 FreeSans 448 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 172816 0 172928 800 0 FreeSans 448 90 0 0 irq[0]
port 114 nsew signal tristate
flabel metal2 s 173376 0 173488 800 0 FreeSans 448 90 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 173936 0 174048 800 0 FreeSans 448 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 65296 0 65408 800 0 FreeSans 448 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 82096 0 82208 800 0 FreeSans 448 90 0 0 la_data_in[10]
port 118 nsew signal input
flabel metal2 s 83776 0 83888 800 0 FreeSans 448 90 0 0 la_data_in[11]
port 119 nsew signal input
flabel metal2 s 85456 0 85568 800 0 FreeSans 448 90 0 0 la_data_in[12]
port 120 nsew signal input
flabel metal2 s 87136 0 87248 800 0 FreeSans 448 90 0 0 la_data_in[13]
port 121 nsew signal input
flabel metal2 s 88816 0 88928 800 0 FreeSans 448 90 0 0 la_data_in[14]
port 122 nsew signal input
flabel metal2 s 90496 0 90608 800 0 FreeSans 448 90 0 0 la_data_in[15]
port 123 nsew signal input
flabel metal2 s 92176 0 92288 800 0 FreeSans 448 90 0 0 la_data_in[16]
port 124 nsew signal input
flabel metal2 s 93856 0 93968 800 0 FreeSans 448 90 0 0 la_data_in[17]
port 125 nsew signal input
flabel metal2 s 95536 0 95648 800 0 FreeSans 448 90 0 0 la_data_in[18]
port 126 nsew signal input
flabel metal2 s 97216 0 97328 800 0 FreeSans 448 90 0 0 la_data_in[19]
port 127 nsew signal input
flabel metal2 s 66976 0 67088 800 0 FreeSans 448 90 0 0 la_data_in[1]
port 128 nsew signal input
flabel metal2 s 98896 0 99008 800 0 FreeSans 448 90 0 0 la_data_in[20]
port 129 nsew signal input
flabel metal2 s 100576 0 100688 800 0 FreeSans 448 90 0 0 la_data_in[21]
port 130 nsew signal input
flabel metal2 s 102256 0 102368 800 0 FreeSans 448 90 0 0 la_data_in[22]
port 131 nsew signal input
flabel metal2 s 103936 0 104048 800 0 FreeSans 448 90 0 0 la_data_in[23]
port 132 nsew signal input
flabel metal2 s 105616 0 105728 800 0 FreeSans 448 90 0 0 la_data_in[24]
port 133 nsew signal input
flabel metal2 s 107296 0 107408 800 0 FreeSans 448 90 0 0 la_data_in[25]
port 134 nsew signal input
flabel metal2 s 108976 0 109088 800 0 FreeSans 448 90 0 0 la_data_in[26]
port 135 nsew signal input
flabel metal2 s 110656 0 110768 800 0 FreeSans 448 90 0 0 la_data_in[27]
port 136 nsew signal input
flabel metal2 s 112336 0 112448 800 0 FreeSans 448 90 0 0 la_data_in[28]
port 137 nsew signal input
flabel metal2 s 114016 0 114128 800 0 FreeSans 448 90 0 0 la_data_in[29]
port 138 nsew signal input
flabel metal2 s 68656 0 68768 800 0 FreeSans 448 90 0 0 la_data_in[2]
port 139 nsew signal input
flabel metal2 s 115696 0 115808 800 0 FreeSans 448 90 0 0 la_data_in[30]
port 140 nsew signal input
flabel metal2 s 117376 0 117488 800 0 FreeSans 448 90 0 0 la_data_in[31]
port 141 nsew signal input
flabel metal2 s 119056 0 119168 800 0 FreeSans 448 90 0 0 la_data_in[32]
port 142 nsew signal input
flabel metal2 s 120736 0 120848 800 0 FreeSans 448 90 0 0 la_data_in[33]
port 143 nsew signal input
flabel metal2 s 122416 0 122528 800 0 FreeSans 448 90 0 0 la_data_in[34]
port 144 nsew signal input
flabel metal2 s 124096 0 124208 800 0 FreeSans 448 90 0 0 la_data_in[35]
port 145 nsew signal input
flabel metal2 s 125776 0 125888 800 0 FreeSans 448 90 0 0 la_data_in[36]
port 146 nsew signal input
flabel metal2 s 127456 0 127568 800 0 FreeSans 448 90 0 0 la_data_in[37]
port 147 nsew signal input
flabel metal2 s 129136 0 129248 800 0 FreeSans 448 90 0 0 la_data_in[38]
port 148 nsew signal input
flabel metal2 s 130816 0 130928 800 0 FreeSans 448 90 0 0 la_data_in[39]
port 149 nsew signal input
flabel metal2 s 70336 0 70448 800 0 FreeSans 448 90 0 0 la_data_in[3]
port 150 nsew signal input
flabel metal2 s 132496 0 132608 800 0 FreeSans 448 90 0 0 la_data_in[40]
port 151 nsew signal input
flabel metal2 s 134176 0 134288 800 0 FreeSans 448 90 0 0 la_data_in[41]
port 152 nsew signal input
flabel metal2 s 135856 0 135968 800 0 FreeSans 448 90 0 0 la_data_in[42]
port 153 nsew signal input
flabel metal2 s 137536 0 137648 800 0 FreeSans 448 90 0 0 la_data_in[43]
port 154 nsew signal input
flabel metal2 s 139216 0 139328 800 0 FreeSans 448 90 0 0 la_data_in[44]
port 155 nsew signal input
flabel metal2 s 140896 0 141008 800 0 FreeSans 448 90 0 0 la_data_in[45]
port 156 nsew signal input
flabel metal2 s 142576 0 142688 800 0 FreeSans 448 90 0 0 la_data_in[46]
port 157 nsew signal input
flabel metal2 s 144256 0 144368 800 0 FreeSans 448 90 0 0 la_data_in[47]
port 158 nsew signal input
flabel metal2 s 145936 0 146048 800 0 FreeSans 448 90 0 0 la_data_in[48]
port 159 nsew signal input
flabel metal2 s 147616 0 147728 800 0 FreeSans 448 90 0 0 la_data_in[49]
port 160 nsew signal input
flabel metal2 s 72016 0 72128 800 0 FreeSans 448 90 0 0 la_data_in[4]
port 161 nsew signal input
flabel metal2 s 149296 0 149408 800 0 FreeSans 448 90 0 0 la_data_in[50]
port 162 nsew signal input
flabel metal2 s 150976 0 151088 800 0 FreeSans 448 90 0 0 la_data_in[51]
port 163 nsew signal input
flabel metal2 s 152656 0 152768 800 0 FreeSans 448 90 0 0 la_data_in[52]
port 164 nsew signal input
flabel metal2 s 154336 0 154448 800 0 FreeSans 448 90 0 0 la_data_in[53]
port 165 nsew signal input
flabel metal2 s 156016 0 156128 800 0 FreeSans 448 90 0 0 la_data_in[54]
port 166 nsew signal input
flabel metal2 s 157696 0 157808 800 0 FreeSans 448 90 0 0 la_data_in[55]
port 167 nsew signal input
flabel metal2 s 159376 0 159488 800 0 FreeSans 448 90 0 0 la_data_in[56]
port 168 nsew signal input
flabel metal2 s 161056 0 161168 800 0 FreeSans 448 90 0 0 la_data_in[57]
port 169 nsew signal input
flabel metal2 s 162736 0 162848 800 0 FreeSans 448 90 0 0 la_data_in[58]
port 170 nsew signal input
flabel metal2 s 164416 0 164528 800 0 FreeSans 448 90 0 0 la_data_in[59]
port 171 nsew signal input
flabel metal2 s 73696 0 73808 800 0 FreeSans 448 90 0 0 la_data_in[5]
port 172 nsew signal input
flabel metal2 s 166096 0 166208 800 0 FreeSans 448 90 0 0 la_data_in[60]
port 173 nsew signal input
flabel metal2 s 167776 0 167888 800 0 FreeSans 448 90 0 0 la_data_in[61]
port 174 nsew signal input
flabel metal2 s 169456 0 169568 800 0 FreeSans 448 90 0 0 la_data_in[62]
port 175 nsew signal input
flabel metal2 s 171136 0 171248 800 0 FreeSans 448 90 0 0 la_data_in[63]
port 176 nsew signal input
flabel metal2 s 75376 0 75488 800 0 FreeSans 448 90 0 0 la_data_in[6]
port 177 nsew signal input
flabel metal2 s 77056 0 77168 800 0 FreeSans 448 90 0 0 la_data_in[7]
port 178 nsew signal input
flabel metal2 s 78736 0 78848 800 0 FreeSans 448 90 0 0 la_data_in[8]
port 179 nsew signal input
flabel metal2 s 80416 0 80528 800 0 FreeSans 448 90 0 0 la_data_in[9]
port 180 nsew signal input
flabel metal2 s 65856 0 65968 800 0 FreeSans 448 90 0 0 la_data_out[0]
port 181 nsew signal tristate
flabel metal2 s 82656 0 82768 800 0 FreeSans 448 90 0 0 la_data_out[10]
port 182 nsew signal tristate
flabel metal2 s 84336 0 84448 800 0 FreeSans 448 90 0 0 la_data_out[11]
port 183 nsew signal tristate
flabel metal2 s 86016 0 86128 800 0 FreeSans 448 90 0 0 la_data_out[12]
port 184 nsew signal tristate
flabel metal2 s 87696 0 87808 800 0 FreeSans 448 90 0 0 la_data_out[13]
port 185 nsew signal tristate
flabel metal2 s 89376 0 89488 800 0 FreeSans 448 90 0 0 la_data_out[14]
port 186 nsew signal tristate
flabel metal2 s 91056 0 91168 800 0 FreeSans 448 90 0 0 la_data_out[15]
port 187 nsew signal tristate
flabel metal2 s 92736 0 92848 800 0 FreeSans 448 90 0 0 la_data_out[16]
port 188 nsew signal tristate
flabel metal2 s 94416 0 94528 800 0 FreeSans 448 90 0 0 la_data_out[17]
port 189 nsew signal tristate
flabel metal2 s 96096 0 96208 800 0 FreeSans 448 90 0 0 la_data_out[18]
port 190 nsew signal tristate
flabel metal2 s 97776 0 97888 800 0 FreeSans 448 90 0 0 la_data_out[19]
port 191 nsew signal tristate
flabel metal2 s 67536 0 67648 800 0 FreeSans 448 90 0 0 la_data_out[1]
port 192 nsew signal tristate
flabel metal2 s 99456 0 99568 800 0 FreeSans 448 90 0 0 la_data_out[20]
port 193 nsew signal tristate
flabel metal2 s 101136 0 101248 800 0 FreeSans 448 90 0 0 la_data_out[21]
port 194 nsew signal tristate
flabel metal2 s 102816 0 102928 800 0 FreeSans 448 90 0 0 la_data_out[22]
port 195 nsew signal tristate
flabel metal2 s 104496 0 104608 800 0 FreeSans 448 90 0 0 la_data_out[23]
port 196 nsew signal tristate
flabel metal2 s 106176 0 106288 800 0 FreeSans 448 90 0 0 la_data_out[24]
port 197 nsew signal tristate
flabel metal2 s 107856 0 107968 800 0 FreeSans 448 90 0 0 la_data_out[25]
port 198 nsew signal tristate
flabel metal2 s 109536 0 109648 800 0 FreeSans 448 90 0 0 la_data_out[26]
port 199 nsew signal tristate
flabel metal2 s 111216 0 111328 800 0 FreeSans 448 90 0 0 la_data_out[27]
port 200 nsew signal tristate
flabel metal2 s 112896 0 113008 800 0 FreeSans 448 90 0 0 la_data_out[28]
port 201 nsew signal tristate
flabel metal2 s 114576 0 114688 800 0 FreeSans 448 90 0 0 la_data_out[29]
port 202 nsew signal tristate
flabel metal2 s 69216 0 69328 800 0 FreeSans 448 90 0 0 la_data_out[2]
port 203 nsew signal tristate
flabel metal2 s 116256 0 116368 800 0 FreeSans 448 90 0 0 la_data_out[30]
port 204 nsew signal tristate
flabel metal2 s 117936 0 118048 800 0 FreeSans 448 90 0 0 la_data_out[31]
port 205 nsew signal tristate
flabel metal2 s 119616 0 119728 800 0 FreeSans 448 90 0 0 la_data_out[32]
port 206 nsew signal tristate
flabel metal2 s 121296 0 121408 800 0 FreeSans 448 90 0 0 la_data_out[33]
port 207 nsew signal tristate
flabel metal2 s 122976 0 123088 800 0 FreeSans 448 90 0 0 la_data_out[34]
port 208 nsew signal tristate
flabel metal2 s 124656 0 124768 800 0 FreeSans 448 90 0 0 la_data_out[35]
port 209 nsew signal tristate
flabel metal2 s 126336 0 126448 800 0 FreeSans 448 90 0 0 la_data_out[36]
port 210 nsew signal tristate
flabel metal2 s 128016 0 128128 800 0 FreeSans 448 90 0 0 la_data_out[37]
port 211 nsew signal tristate
flabel metal2 s 129696 0 129808 800 0 FreeSans 448 90 0 0 la_data_out[38]
port 212 nsew signal tristate
flabel metal2 s 131376 0 131488 800 0 FreeSans 448 90 0 0 la_data_out[39]
port 213 nsew signal tristate
flabel metal2 s 70896 0 71008 800 0 FreeSans 448 90 0 0 la_data_out[3]
port 214 nsew signal tristate
flabel metal2 s 133056 0 133168 800 0 FreeSans 448 90 0 0 la_data_out[40]
port 215 nsew signal tristate
flabel metal2 s 134736 0 134848 800 0 FreeSans 448 90 0 0 la_data_out[41]
port 216 nsew signal tristate
flabel metal2 s 136416 0 136528 800 0 FreeSans 448 90 0 0 la_data_out[42]
port 217 nsew signal tristate
flabel metal2 s 138096 0 138208 800 0 FreeSans 448 90 0 0 la_data_out[43]
port 218 nsew signal tristate
flabel metal2 s 139776 0 139888 800 0 FreeSans 448 90 0 0 la_data_out[44]
port 219 nsew signal tristate
flabel metal2 s 141456 0 141568 800 0 FreeSans 448 90 0 0 la_data_out[45]
port 220 nsew signal tristate
flabel metal2 s 143136 0 143248 800 0 FreeSans 448 90 0 0 la_data_out[46]
port 221 nsew signal tristate
flabel metal2 s 144816 0 144928 800 0 FreeSans 448 90 0 0 la_data_out[47]
port 222 nsew signal tristate
flabel metal2 s 146496 0 146608 800 0 FreeSans 448 90 0 0 la_data_out[48]
port 223 nsew signal tristate
flabel metal2 s 148176 0 148288 800 0 FreeSans 448 90 0 0 la_data_out[49]
port 224 nsew signal tristate
flabel metal2 s 72576 0 72688 800 0 FreeSans 448 90 0 0 la_data_out[4]
port 225 nsew signal tristate
flabel metal2 s 149856 0 149968 800 0 FreeSans 448 90 0 0 la_data_out[50]
port 226 nsew signal tristate
flabel metal2 s 151536 0 151648 800 0 FreeSans 448 90 0 0 la_data_out[51]
port 227 nsew signal tristate
flabel metal2 s 153216 0 153328 800 0 FreeSans 448 90 0 0 la_data_out[52]
port 228 nsew signal tristate
flabel metal2 s 154896 0 155008 800 0 FreeSans 448 90 0 0 la_data_out[53]
port 229 nsew signal tristate
flabel metal2 s 156576 0 156688 800 0 FreeSans 448 90 0 0 la_data_out[54]
port 230 nsew signal tristate
flabel metal2 s 158256 0 158368 800 0 FreeSans 448 90 0 0 la_data_out[55]
port 231 nsew signal tristate
flabel metal2 s 159936 0 160048 800 0 FreeSans 448 90 0 0 la_data_out[56]
port 232 nsew signal tristate
flabel metal2 s 161616 0 161728 800 0 FreeSans 448 90 0 0 la_data_out[57]
port 233 nsew signal tristate
flabel metal2 s 163296 0 163408 800 0 FreeSans 448 90 0 0 la_data_out[58]
port 234 nsew signal tristate
flabel metal2 s 164976 0 165088 800 0 FreeSans 448 90 0 0 la_data_out[59]
port 235 nsew signal tristate
flabel metal2 s 74256 0 74368 800 0 FreeSans 448 90 0 0 la_data_out[5]
port 236 nsew signal tristate
flabel metal2 s 166656 0 166768 800 0 FreeSans 448 90 0 0 la_data_out[60]
port 237 nsew signal tristate
flabel metal2 s 168336 0 168448 800 0 FreeSans 448 90 0 0 la_data_out[61]
port 238 nsew signal tristate
flabel metal2 s 170016 0 170128 800 0 FreeSans 448 90 0 0 la_data_out[62]
port 239 nsew signal tristate
flabel metal2 s 171696 0 171808 800 0 FreeSans 448 90 0 0 la_data_out[63]
port 240 nsew signal tristate
flabel metal2 s 75936 0 76048 800 0 FreeSans 448 90 0 0 la_data_out[6]
port 241 nsew signal tristate
flabel metal2 s 77616 0 77728 800 0 FreeSans 448 90 0 0 la_data_out[7]
port 242 nsew signal tristate
flabel metal2 s 79296 0 79408 800 0 FreeSans 448 90 0 0 la_data_out[8]
port 243 nsew signal tristate
flabel metal2 s 80976 0 81088 800 0 FreeSans 448 90 0 0 la_data_out[9]
port 244 nsew signal tristate
flabel metal2 s 66416 0 66528 800 0 FreeSans 448 90 0 0 la_oenb[0]
port 245 nsew signal input
flabel metal2 s 83216 0 83328 800 0 FreeSans 448 90 0 0 la_oenb[10]
port 246 nsew signal input
flabel metal2 s 84896 0 85008 800 0 FreeSans 448 90 0 0 la_oenb[11]
port 247 nsew signal input
flabel metal2 s 86576 0 86688 800 0 FreeSans 448 90 0 0 la_oenb[12]
port 248 nsew signal input
flabel metal2 s 88256 0 88368 800 0 FreeSans 448 90 0 0 la_oenb[13]
port 249 nsew signal input
flabel metal2 s 89936 0 90048 800 0 FreeSans 448 90 0 0 la_oenb[14]
port 250 nsew signal input
flabel metal2 s 91616 0 91728 800 0 FreeSans 448 90 0 0 la_oenb[15]
port 251 nsew signal input
flabel metal2 s 93296 0 93408 800 0 FreeSans 448 90 0 0 la_oenb[16]
port 252 nsew signal input
flabel metal2 s 94976 0 95088 800 0 FreeSans 448 90 0 0 la_oenb[17]
port 253 nsew signal input
flabel metal2 s 96656 0 96768 800 0 FreeSans 448 90 0 0 la_oenb[18]
port 254 nsew signal input
flabel metal2 s 98336 0 98448 800 0 FreeSans 448 90 0 0 la_oenb[19]
port 255 nsew signal input
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 la_oenb[1]
port 256 nsew signal input
flabel metal2 s 100016 0 100128 800 0 FreeSans 448 90 0 0 la_oenb[20]
port 257 nsew signal input
flabel metal2 s 101696 0 101808 800 0 FreeSans 448 90 0 0 la_oenb[21]
port 258 nsew signal input
flabel metal2 s 103376 0 103488 800 0 FreeSans 448 90 0 0 la_oenb[22]
port 259 nsew signal input
flabel metal2 s 105056 0 105168 800 0 FreeSans 448 90 0 0 la_oenb[23]
port 260 nsew signal input
flabel metal2 s 106736 0 106848 800 0 FreeSans 448 90 0 0 la_oenb[24]
port 261 nsew signal input
flabel metal2 s 108416 0 108528 800 0 FreeSans 448 90 0 0 la_oenb[25]
port 262 nsew signal input
flabel metal2 s 110096 0 110208 800 0 FreeSans 448 90 0 0 la_oenb[26]
port 263 nsew signal input
flabel metal2 s 111776 0 111888 800 0 FreeSans 448 90 0 0 la_oenb[27]
port 264 nsew signal input
flabel metal2 s 113456 0 113568 800 0 FreeSans 448 90 0 0 la_oenb[28]
port 265 nsew signal input
flabel metal2 s 115136 0 115248 800 0 FreeSans 448 90 0 0 la_oenb[29]
port 266 nsew signal input
flabel metal2 s 69776 0 69888 800 0 FreeSans 448 90 0 0 la_oenb[2]
port 267 nsew signal input
flabel metal2 s 116816 0 116928 800 0 FreeSans 448 90 0 0 la_oenb[30]
port 268 nsew signal input
flabel metal2 s 118496 0 118608 800 0 FreeSans 448 90 0 0 la_oenb[31]
port 269 nsew signal input
flabel metal2 s 120176 0 120288 800 0 FreeSans 448 90 0 0 la_oenb[32]
port 270 nsew signal input
flabel metal2 s 121856 0 121968 800 0 FreeSans 448 90 0 0 la_oenb[33]
port 271 nsew signal input
flabel metal2 s 123536 0 123648 800 0 FreeSans 448 90 0 0 la_oenb[34]
port 272 nsew signal input
flabel metal2 s 125216 0 125328 800 0 FreeSans 448 90 0 0 la_oenb[35]
port 273 nsew signal input
flabel metal2 s 126896 0 127008 800 0 FreeSans 448 90 0 0 la_oenb[36]
port 274 nsew signal input
flabel metal2 s 128576 0 128688 800 0 FreeSans 448 90 0 0 la_oenb[37]
port 275 nsew signal input
flabel metal2 s 130256 0 130368 800 0 FreeSans 448 90 0 0 la_oenb[38]
port 276 nsew signal input
flabel metal2 s 131936 0 132048 800 0 FreeSans 448 90 0 0 la_oenb[39]
port 277 nsew signal input
flabel metal2 s 71456 0 71568 800 0 FreeSans 448 90 0 0 la_oenb[3]
port 278 nsew signal input
flabel metal2 s 133616 0 133728 800 0 FreeSans 448 90 0 0 la_oenb[40]
port 279 nsew signal input
flabel metal2 s 135296 0 135408 800 0 FreeSans 448 90 0 0 la_oenb[41]
port 280 nsew signal input
flabel metal2 s 136976 0 137088 800 0 FreeSans 448 90 0 0 la_oenb[42]
port 281 nsew signal input
flabel metal2 s 138656 0 138768 800 0 FreeSans 448 90 0 0 la_oenb[43]
port 282 nsew signal input
flabel metal2 s 140336 0 140448 800 0 FreeSans 448 90 0 0 la_oenb[44]
port 283 nsew signal input
flabel metal2 s 142016 0 142128 800 0 FreeSans 448 90 0 0 la_oenb[45]
port 284 nsew signal input
flabel metal2 s 143696 0 143808 800 0 FreeSans 448 90 0 0 la_oenb[46]
port 285 nsew signal input
flabel metal2 s 145376 0 145488 800 0 FreeSans 448 90 0 0 la_oenb[47]
port 286 nsew signal input
flabel metal2 s 147056 0 147168 800 0 FreeSans 448 90 0 0 la_oenb[48]
port 287 nsew signal input
flabel metal2 s 148736 0 148848 800 0 FreeSans 448 90 0 0 la_oenb[49]
port 288 nsew signal input
flabel metal2 s 73136 0 73248 800 0 FreeSans 448 90 0 0 la_oenb[4]
port 289 nsew signal input
flabel metal2 s 150416 0 150528 800 0 FreeSans 448 90 0 0 la_oenb[50]
port 290 nsew signal input
flabel metal2 s 152096 0 152208 800 0 FreeSans 448 90 0 0 la_oenb[51]
port 291 nsew signal input
flabel metal2 s 153776 0 153888 800 0 FreeSans 448 90 0 0 la_oenb[52]
port 292 nsew signal input
flabel metal2 s 155456 0 155568 800 0 FreeSans 448 90 0 0 la_oenb[53]
port 293 nsew signal input
flabel metal2 s 157136 0 157248 800 0 FreeSans 448 90 0 0 la_oenb[54]
port 294 nsew signal input
flabel metal2 s 158816 0 158928 800 0 FreeSans 448 90 0 0 la_oenb[55]
port 295 nsew signal input
flabel metal2 s 160496 0 160608 800 0 FreeSans 448 90 0 0 la_oenb[56]
port 296 nsew signal input
flabel metal2 s 162176 0 162288 800 0 FreeSans 448 90 0 0 la_oenb[57]
port 297 nsew signal input
flabel metal2 s 163856 0 163968 800 0 FreeSans 448 90 0 0 la_oenb[58]
port 298 nsew signal input
flabel metal2 s 165536 0 165648 800 0 FreeSans 448 90 0 0 la_oenb[59]
port 299 nsew signal input
flabel metal2 s 74816 0 74928 800 0 FreeSans 448 90 0 0 la_oenb[5]
port 300 nsew signal input
flabel metal2 s 167216 0 167328 800 0 FreeSans 448 90 0 0 la_oenb[60]
port 301 nsew signal input
flabel metal2 s 168896 0 169008 800 0 FreeSans 448 90 0 0 la_oenb[61]
port 302 nsew signal input
flabel metal2 s 170576 0 170688 800 0 FreeSans 448 90 0 0 la_oenb[62]
port 303 nsew signal input
flabel metal2 s 172256 0 172368 800 0 FreeSans 448 90 0 0 la_oenb[63]
port 304 nsew signal input
flabel metal2 s 76496 0 76608 800 0 FreeSans 448 90 0 0 la_oenb[6]
port 305 nsew signal input
flabel metal2 s 78176 0 78288 800 0 FreeSans 448 90 0 0 la_oenb[7]
port 306 nsew signal input
flabel metal2 s 79856 0 79968 800 0 FreeSans 448 90 0 0 la_oenb[8]
port 307 nsew signal input
flabel metal2 s 81536 0 81648 800 0 FreeSans 448 90 0 0 la_oenb[9]
port 308 nsew signal input
flabel metal4 s 4448 3076 4768 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 35168 3076 35488 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 65888 3076 66208 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 96608 3076 96928 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 127328 3076 127648 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 158048 3076 158368 116876 0 FreeSans 1280 90 0 0 vdd
port 309 nsew power bidirectional
flabel metal4 s 19808 3076 20128 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 81248 3076 81568 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 111968 3076 112288 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 142688 3076 143008 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal4 s 173408 3076 173728 116876 0 FreeSans 1280 90 0 0 vss
port 310 nsew ground bidirectional
flabel metal2 s 5936 0 6048 800 0 FreeSans 448 90 0 0 wb_clk_i
port 311 nsew signal input
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 wb_rst_i
port 312 nsew signal input
flabel metal2 s 7056 0 7168 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 313 nsew signal tristate
flabel metal2 s 9296 0 9408 800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 314 nsew signal input
flabel metal2 s 28336 0 28448 800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 315 nsew signal input
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 316 nsew signal input
flabel metal2 s 31696 0 31808 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 317 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 318 nsew signal input
flabel metal2 s 35056 0 35168 800 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 319 nsew signal input
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 320 nsew signal input
flabel metal2 s 38416 0 38528 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 321 nsew signal input
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 322 nsew signal input
flabel metal2 s 41776 0 41888 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 323 nsew signal input
flabel metal2 s 43456 0 43568 800 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 324 nsew signal input
flabel metal2 s 11536 0 11648 800 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 325 nsew signal input
flabel metal2 s 45136 0 45248 800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 326 nsew signal input
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 327 nsew signal input
flabel metal2 s 48496 0 48608 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 328 nsew signal input
flabel metal2 s 50176 0 50288 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 329 nsew signal input
flabel metal2 s 51856 0 51968 800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 330 nsew signal input
flabel metal2 s 53536 0 53648 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 331 nsew signal input
flabel metal2 s 55216 0 55328 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 332 nsew signal input
flabel metal2 s 56896 0 57008 800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 333 nsew signal input
flabel metal2 s 58576 0 58688 800 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 334 nsew signal input
flabel metal2 s 60256 0 60368 800 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 335 nsew signal input
flabel metal2 s 13776 0 13888 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 336 nsew signal input
flabel metal2 s 61936 0 62048 800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 337 nsew signal input
flabel metal2 s 63616 0 63728 800 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 338 nsew signal input
flabel metal2 s 16016 0 16128 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 339 nsew signal input
flabel metal2 s 18256 0 18368 800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 340 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 341 nsew signal input
flabel metal2 s 21616 0 21728 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 342 nsew signal input
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 343 nsew signal input
flabel metal2 s 24976 0 25088 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 344 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 345 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 346 nsew signal input
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 347 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 348 nsew signal input
flabel metal2 s 30576 0 30688 800 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 349 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 350 nsew signal input
flabel metal2 s 33936 0 34048 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 351 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 352 nsew signal input
flabel metal2 s 37296 0 37408 800 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 353 nsew signal input
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 354 nsew signal input
flabel metal2 s 40656 0 40768 800 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 355 nsew signal input
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 356 nsew signal input
flabel metal2 s 44016 0 44128 800 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 357 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 358 nsew signal input
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 359 nsew signal input
flabel metal2 s 47376 0 47488 800 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 360 nsew signal input
flabel metal2 s 49056 0 49168 800 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 361 nsew signal input
flabel metal2 s 50736 0 50848 800 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 362 nsew signal input
flabel metal2 s 52416 0 52528 800 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 363 nsew signal input
flabel metal2 s 54096 0 54208 800 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 364 nsew signal input
flabel metal2 s 55776 0 55888 800 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 365 nsew signal input
flabel metal2 s 57456 0 57568 800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 366 nsew signal input
flabel metal2 s 59136 0 59248 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 367 nsew signal input
flabel metal2 s 60816 0 60928 800 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 368 nsew signal input
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 369 nsew signal input
flabel metal2 s 62496 0 62608 800 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 370 nsew signal input
flabel metal2 s 64176 0 64288 800 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 371 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 372 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 373 nsew signal input
flabel metal2 s 20496 0 20608 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 374 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 375 nsew signal input
flabel metal2 s 23856 0 23968 800 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 376 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 377 nsew signal input
flabel metal2 s 27216 0 27328 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 378 nsew signal input
flabel metal2 s 10416 0 10528 800 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 379 nsew signal tristate
flabel metal2 s 29456 0 29568 800 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 380 nsew signal tristate
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 381 nsew signal tristate
flabel metal2 s 32816 0 32928 800 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 382 nsew signal tristate
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 383 nsew signal tristate
flabel metal2 s 36176 0 36288 800 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 384 nsew signal tristate
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 385 nsew signal tristate
flabel metal2 s 39536 0 39648 800 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 386 nsew signal tristate
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 387 nsew signal tristate
flabel metal2 s 42896 0 43008 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 388 nsew signal tristate
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 389 nsew signal tristate
flabel metal2 s 12656 0 12768 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 390 nsew signal tristate
flabel metal2 s 46256 0 46368 800 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 391 nsew signal tristate
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 392 nsew signal tristate
flabel metal2 s 49616 0 49728 800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 393 nsew signal tristate
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 394 nsew signal tristate
flabel metal2 s 52976 0 53088 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 395 nsew signal tristate
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 396 nsew signal tristate
flabel metal2 s 56336 0 56448 800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 397 nsew signal tristate
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 398 nsew signal tristate
flabel metal2 s 59696 0 59808 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 399 nsew signal tristate
flabel metal2 s 61376 0 61488 800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 400 nsew signal tristate
flabel metal2 s 14896 0 15008 800 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 401 nsew signal tristate
flabel metal2 s 63056 0 63168 800 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 402 nsew signal tristate
flabel metal2 s 64736 0 64848 800 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 403 nsew signal tristate
flabel metal2 s 17136 0 17248 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 404 nsew signal tristate
flabel metal2 s 19376 0 19488 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 405 nsew signal tristate
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 406 nsew signal tristate
flabel metal2 s 22736 0 22848 800 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 407 nsew signal tristate
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 408 nsew signal tristate
flabel metal2 s 26096 0 26208 800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 409 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 410 nsew signal tristate
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 411 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 412 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 413 nsew signal input
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 414 nsew signal input
flabel metal2 s 8176 0 8288 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 415 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 wbs_we_i
port 416 nsew signal input
rlabel metal1 89992 116816 89992 116816 0 vdd
rlabel metal1 89992 116032 89992 116032 0 vss
rlabel metal3 36960 6664 36960 6664 0 _000_
rlabel metal3 59024 5208 59024 5208 0 _001_
rlabel metal2 66808 9296 66808 9296 0 _002_
rlabel metal3 68152 8904 68152 8904 0 _003_
rlabel metal2 67928 9856 67928 9856 0 _004_
rlabel metal2 71792 9128 71792 9128 0 _005_
rlabel metal2 71848 10304 71848 10304 0 _006_
rlabel metal2 73640 10136 73640 10136 0 _007_
rlabel metal2 76160 9128 76160 9128 0 _008_
rlabel metal2 78680 10024 78680 10024 0 _009_
rlabel metal2 85736 8624 85736 8624 0 _010_
rlabel metal3 82656 10024 82656 10024 0 _011_
rlabel metal2 86408 10864 86408 10864 0 _012_
rlabel metal3 88368 9688 88368 9688 0 _013_
rlabel metal3 89992 10472 89992 10472 0 _014_
rlabel metal2 83552 10696 83552 10696 0 _015_
rlabel metal2 91560 11480 91560 11480 0 _016_
rlabel metal2 104328 11032 104328 11032 0 _017_
rlabel metal2 105448 11424 105448 11424 0 _018_
rlabel metal2 112728 11088 112728 11088 0 _019_
rlabel metal3 115752 9576 115752 9576 0 _020_
rlabel metal2 113176 10360 113176 10360 0 _021_
rlabel metal2 115864 8288 115864 8288 0 _022_
rlabel metal3 114688 12040 114688 12040 0 _023_
rlabel metal2 110264 5544 110264 5544 0 _024_
rlabel metal2 109368 7000 109368 7000 0 _025_
rlabel metal2 103432 8288 103432 8288 0 _026_
rlabel metal2 105224 8456 105224 8456 0 _027_
rlabel metal2 95480 10416 95480 10416 0 _028_
rlabel metal2 91896 8456 91896 8456 0 _029_
rlabel metal2 99288 11760 99288 11760 0 _030_
rlabel metal2 101864 9520 101864 9520 0 _031_
rlabel metal2 99792 9240 99792 9240 0 _032_
rlabel metal3 36624 4984 36624 4984 0 _033_
rlabel metal3 60144 4424 60144 4424 0 _034_
rlabel metal2 12824 4648 12824 4648 0 _035_
rlabel metal2 16632 4816 16632 4816 0 _036_
rlabel metal2 18984 7784 18984 7784 0 _037_
rlabel metal2 20216 5264 20216 5264 0 _038_
rlabel metal2 26488 6216 26488 6216 0 _039_
rlabel metal2 37800 6216 37800 6216 0 _040_
rlabel metal2 26040 4760 26040 4760 0 _041_
rlabel metal2 26488 7784 26488 7784 0 _042_
rlabel metal3 35224 6552 35224 6552 0 _043_
rlabel metal2 29960 4648 29960 4648 0 _044_
rlabel metal2 31864 9464 31864 9464 0 _045_
rlabel metal2 31976 7896 31976 7896 0 _046_
rlabel metal2 45080 5488 45080 5488 0 _047_
rlabel metal2 51240 4480 51240 4480 0 _048_
rlabel metal2 38360 10304 38360 10304 0 _049_
rlabel metal3 38976 8904 38976 8904 0 _050_
rlabel metal3 43512 7560 43512 7560 0 _051_
rlabel metal2 43708 9688 43708 9688 0 _052_
rlabel metal2 50344 8372 50344 8372 0 _053_
rlabel metal2 47432 10304 47432 10304 0 _054_
rlabel metal2 47712 4424 47712 4424 0 _055_
rlabel metal2 51912 6608 51912 6608 0 _056_
rlabel metal2 53256 10920 53256 10920 0 _057_
rlabel metal2 57960 5488 57960 5488 0 _058_
rlabel metal2 54264 7336 54264 7336 0 _059_
rlabel metal2 56952 10304 56952 10304 0 _060_
rlabel metal2 60536 10136 60536 10136 0 _061_
rlabel metal2 61656 6216 61656 6216 0 _062_
rlabel metal3 61880 7672 61880 7672 0 _063_
rlabel metal2 63000 6888 63000 6888 0 _064_
rlabel metal3 91112 4312 91112 4312 0 _065_
rlabel metal2 140952 5544 140952 5544 0 _066_
rlabel metal2 133896 4592 133896 4592 0 _067_
rlabel metal3 133896 6384 133896 6384 0 _068_
rlabel metal2 137368 7168 137368 7168 0 _069_
rlabel metal3 70616 4312 70616 4312 0 _070_
rlabel metal3 49560 6552 49560 6552 0 _071_
rlabel metal2 48104 6328 48104 6328 0 _072_
rlabel metal2 44856 9072 44856 9072 0 _073_
rlabel metal2 116088 10136 116088 10136 0 _074_
rlabel metal2 59472 6104 59472 6104 0 _075_
rlabel metal3 68320 6104 68320 6104 0 _076_
rlabel metal3 128800 5880 128800 5880 0 _077_
rlabel metal3 127456 4424 127456 4424 0 _078_
rlabel metal2 125048 6440 125048 6440 0 _079_
rlabel metal2 70112 5208 70112 5208 0 _080_
rlabel metal2 124040 5040 124040 5040 0 _081_
rlabel metal2 123592 4144 123592 4144 0 _082_
rlabel metal3 143304 4984 143304 4984 0 _083_
rlabel metal2 141736 6328 141736 6328 0 _084_
rlabel metal3 103040 2744 103040 2744 0 _085_
rlabel metal2 68152 4480 68152 4480 0 _086_
rlabel metal3 115808 6104 115808 6104 0 _087_
rlabel metal3 106008 20664 106008 20664 0 _088_
rlabel metal2 139272 3864 139272 3864 0 _089_
rlabel metal3 106344 19208 106344 19208 0 _090_
rlabel metal2 101640 11032 101640 11032 0 _091_
rlabel metal2 113064 5880 113064 5880 0 _092_
rlabel metal2 130088 3248 130088 3248 0 _093_
rlabel metal3 129192 4984 129192 4984 0 _094_
rlabel metal3 126336 5096 126336 5096 0 _095_
rlabel metal3 124320 5096 124320 5096 0 _096_
rlabel metal2 138712 6272 138712 6272 0 _097_
rlabel metal3 135352 6664 135352 6664 0 _098_
rlabel metal2 139776 5656 139776 5656 0 _099_
rlabel metal3 111944 17752 111944 17752 0 _100_
rlabel metal2 92008 7280 92008 7280 0 _101_
rlabel metal3 137648 4984 137648 4984 0 _102_
rlabel metal2 138824 4592 138824 4592 0 _103_
rlabel metal2 143976 7168 143976 7168 0 _104_
rlabel metal3 143640 4088 143640 4088 0 _105_
rlabel metal2 141288 6720 141288 6720 0 _106_
rlabel metal3 143024 5320 143024 5320 0 _107_
rlabel metal2 138152 7336 138152 7336 0 _108_
rlabel metal2 138208 4536 138208 4536 0 _109_
rlabel metal2 148344 3304 148344 3304 0 _110_
rlabel metal2 69104 5880 69104 5880 0 _111_
rlabel metal2 147336 3360 147336 3360 0 _112_
rlabel metal3 134008 7672 134008 7672 0 _113_
rlabel metal3 138376 4928 138376 4928 0 _114_
rlabel metal3 142688 4200 142688 4200 0 _115_
rlabel metal3 143080 5096 143080 5096 0 _116_
rlabel metal3 143472 4312 143472 4312 0 _117_
rlabel metal2 141624 4536 141624 4536 0 _118_
rlabel metal3 140168 4536 140168 4536 0 _119_
rlabel metal3 127736 5320 127736 5320 0 _120_
rlabel metal3 102704 22232 102704 22232 0 _121_
rlabel metal2 92008 4424 92008 4424 0 _122_
rlabel metal2 18872 6384 18872 6384 0 _123_
rlabel metal2 39704 4144 39704 4144 0 _124_
rlabel metal3 76496 7448 76496 7448 0 _125_
rlabel metal2 73752 5096 73752 5096 0 _126_
rlabel metal2 71736 4760 71736 4760 0 _127_
rlabel metal2 66808 6216 66808 6216 0 _128_
rlabel metal2 67256 6048 67256 6048 0 _129_
rlabel metal3 63616 5880 63616 5880 0 _130_
rlabel metal2 42392 6272 42392 6272 0 _131_
rlabel metal2 40768 5992 40768 5992 0 _132_
rlabel metal2 58968 5208 58968 5208 0 _133_
rlabel metal2 73752 10192 73752 10192 0 _134_
rlabel metal3 72464 11144 72464 11144 0 _135_
rlabel metal2 67928 6216 67928 6216 0 _136_
rlabel metal2 67368 4648 67368 4648 0 _137_
rlabel metal2 42840 4984 42840 4984 0 _138_
rlabel metal2 67928 4368 67928 4368 0 _139_
rlabel metal2 67816 4704 67816 4704 0 _140_
rlabel metal2 68264 5824 68264 5824 0 _141_
rlabel metal2 74592 9240 74592 9240 0 _142_
rlabel metal3 70392 6272 70392 6272 0 _143_
rlabel metal2 69384 4872 69384 4872 0 _144_
rlabel metal2 69832 6328 69832 6328 0 _145_
rlabel metal3 69328 7224 69328 7224 0 _146_
rlabel metal2 68488 5600 68488 5600 0 _147_
rlabel metal2 69104 5656 69104 5656 0 _148_
rlabel metal2 69496 6608 69496 6608 0 _149_
rlabel metal2 129976 5264 129976 5264 0 _150_
rlabel metal2 72072 5320 72072 5320 0 _151_
rlabel metal2 22008 7280 22008 7280 0 _152_
rlabel metal2 72520 4928 72520 4928 0 _153_
rlabel metal3 71400 4424 71400 4424 0 _154_
rlabel metal3 80696 4984 80696 4984 0 _155_
rlabel metal2 73640 3976 73640 3976 0 _156_
rlabel metal2 72016 11256 72016 11256 0 _157_
rlabel metal2 75432 9408 75432 9408 0 _158_
rlabel metal3 71400 7336 71400 7336 0 _159_
rlabel metal2 72408 6608 72408 6608 0 _160_
rlabel metal2 74760 7896 74760 7896 0 _161_
rlabel metal2 71400 5376 71400 5376 0 _162_
rlabel metal2 72632 5152 72632 5152 0 _163_
rlabel metal2 74200 6664 74200 6664 0 _164_
rlabel metal3 142520 6440 142520 6440 0 _165_
rlabel metal2 68936 4592 68936 4592 0 _166_
rlabel metal2 78904 8624 78904 8624 0 _167_
rlabel metal2 68544 6664 68544 6664 0 _168_
rlabel metal2 76216 5488 76216 5488 0 _169_
rlabel metal3 77560 4984 77560 4984 0 _170_
rlabel metal2 76664 9688 76664 9688 0 _171_
rlabel metal2 15232 6104 15232 6104 0 _172_
rlabel metal3 81424 5880 81424 5880 0 _173_
rlabel metal2 86856 6384 86856 6384 0 _174_
rlabel metal2 86576 6440 86576 6440 0 _175_
rlabel metal2 80696 8288 80696 8288 0 _176_
rlabel metal2 83944 5768 83944 5768 0 _177_
rlabel metal2 85512 5152 85512 5152 0 _178_
rlabel metal3 84840 6440 84840 6440 0 _179_
rlabel metal3 82096 9688 82096 9688 0 _180_
rlabel metal3 81480 8232 81480 8232 0 _181_
rlabel metal2 76552 7672 76552 7672 0 _182_
rlabel metal2 82488 7784 82488 7784 0 _183_
rlabel metal2 84280 8512 84280 8512 0 _184_
rlabel metal3 85120 8232 85120 8232 0 _185_
rlabel metal2 85848 7448 85848 7448 0 _186_
rlabel metal2 86968 8456 86968 8456 0 _187_
rlabel metal2 86184 10024 86184 10024 0 _188_
rlabel metal2 85064 5152 85064 5152 0 _189_
rlabel metal3 84504 4536 84504 4536 0 _190_
rlabel metal2 51632 10360 51632 10360 0 _191_
rlabel metal2 86520 7728 86520 7728 0 _192_
rlabel metal2 87192 6216 87192 6216 0 _193_
rlabel metal3 86240 4872 86240 4872 0 _194_
rlabel metal2 86576 10360 86576 10360 0 _195_
rlabel metal2 89320 8232 89320 8232 0 _196_
rlabel metal2 90440 6664 90440 6664 0 _197_
rlabel metal2 90776 6832 90776 6832 0 _198_
rlabel metal2 90328 8456 90328 8456 0 _199_
rlabel metal2 90664 4648 90664 4648 0 _200_
rlabel metal2 91112 4816 91112 4816 0 _201_
rlabel metal2 91112 11424 91112 11424 0 _202_
rlabel metal2 44968 7448 44968 7448 0 _203_
rlabel metal2 83160 7112 83160 7112 0 _204_
rlabel metal2 88424 6384 88424 6384 0 _205_
rlabel metal2 82824 4368 82824 4368 0 _206_
rlabel metal3 143584 4536 143584 4536 0 _207_
rlabel metal2 143416 5376 143416 5376 0 _208_
rlabel metal2 83720 6104 83720 6104 0 _209_
rlabel metal3 67816 6832 67816 6832 0 _210_
rlabel metal3 90384 4984 90384 4984 0 _211_
rlabel metal2 91448 7392 91448 7392 0 _212_
rlabel metal2 134680 6608 134680 6608 0 _213_
rlabel metal2 16912 6104 16912 6104 0 _214_
rlabel metal3 76776 8232 76776 8232 0 _215_
rlabel metal2 115304 12936 115304 12936 0 _216_
rlabel metal2 117432 5040 117432 5040 0 _217_
rlabel metal2 112616 6216 112616 6216 0 _218_
rlabel metal3 113064 4424 113064 4424 0 _219_
rlabel metal3 96488 20776 96488 20776 0 _220_
rlabel metal2 117544 4704 117544 4704 0 _221_
rlabel metal3 111384 3304 111384 3304 0 _222_
rlabel metal3 118272 5656 118272 5656 0 _223_
rlabel metal2 118552 5376 118552 5376 0 _224_
rlabel metal3 82880 7224 82880 7224 0 _225_
rlabel metal2 91504 4760 91504 4760 0 _226_
rlabel metal2 118776 7728 118776 7728 0 _227_
rlabel metal3 119392 4312 119392 4312 0 _228_
rlabel metal3 114968 9912 114968 9912 0 _229_
rlabel metal3 116984 9688 116984 9688 0 _230_
rlabel metal2 45976 7644 45976 7644 0 _231_
rlabel metal2 121352 6160 121352 6160 0 _232_
rlabel metal2 120904 4704 120904 4704 0 _233_
rlabel metal2 119560 7280 119560 7280 0 _234_
rlabel metal2 120232 7392 120232 7392 0 _235_
rlabel metal3 119280 5880 119280 5880 0 _236_
rlabel metal2 119560 5320 119560 5320 0 _237_
rlabel metal2 118776 8568 118776 8568 0 _238_
rlabel metal3 120904 5040 120904 5040 0 _239_
rlabel metal2 118552 8680 118552 8680 0 _240_
rlabel metal3 117544 6440 117544 6440 0 _241_
rlabel metal3 105112 6552 105112 6552 0 _242_
rlabel metal2 110376 6944 110376 6944 0 _243_
rlabel metal2 115584 6776 115584 6776 0 _244_
rlabel metal2 118888 7784 118888 7784 0 _245_
rlabel metal3 45920 5992 45920 5992 0 _246_
rlabel metal3 115416 4424 115416 4424 0 _247_
rlabel metal2 116872 7112 116872 7112 0 _248_
rlabel metal2 114856 6384 114856 6384 0 _249_
rlabel metal2 142520 9240 142520 9240 0 _250_
rlabel metal2 114968 5264 114968 5264 0 _251_
rlabel metal2 113848 4704 113848 4704 0 _252_
rlabel metal2 113960 4704 113960 4704 0 _253_
rlabel metal2 21672 3416 21672 3416 0 _254_
rlabel metal3 80696 5992 80696 5992 0 _255_
rlabel metal2 93072 7672 93072 7672 0 _256_
rlabel metal2 108584 4816 108584 4816 0 _257_
rlabel metal2 107800 6328 107800 6328 0 _258_
rlabel metal2 108920 4704 108920 4704 0 _259_
rlabel metal2 94696 5376 94696 5376 0 _260_
rlabel metal2 95032 6160 95032 6160 0 _261_
rlabel metal2 109256 4872 109256 4872 0 _262_
rlabel metal3 107296 7672 107296 7672 0 _263_
rlabel metal3 97216 3304 97216 3304 0 _264_
rlabel metal3 58016 5992 58016 5992 0 _265_
rlabel metal2 102088 5712 102088 5712 0 _266_
rlabel metal3 97104 4424 97104 4424 0 _267_
rlabel metal2 52472 12376 52472 12376 0 _268_
rlabel metal2 103096 5320 103096 5320 0 _269_
rlabel metal3 104608 7448 104608 7448 0 _270_
rlabel metal4 95704 8008 95704 8008 0 _271_
rlabel metal2 101752 5712 101752 5712 0 _272_
rlabel metal2 102424 5152 102424 5152 0 _273_
rlabel metal2 56224 5880 56224 5880 0 _274_
rlabel metal2 106008 4928 106008 4928 0 _275_
rlabel metal2 105336 7392 105336 7392 0 _276_
rlabel metal3 60648 9128 60648 9128 0 _277_
rlabel metal2 97384 6328 97384 6328 0 _278_
rlabel metal2 95928 5880 95928 5880 0 _279_
rlabel metal2 96320 5320 96320 5320 0 _280_
rlabel metal2 138880 7672 138880 7672 0 _281_
rlabel metal2 137088 4424 137088 4424 0 _282_
rlabel metal2 96152 6608 96152 6608 0 _283_
rlabel metal3 98168 1624 98168 1624 0 _284_
rlabel metal2 97384 5320 97384 5320 0 _285_
rlabel metal2 93184 8008 93184 8008 0 _286_
rlabel metal2 98840 8736 98840 8736 0 _287_
rlabel metal2 99176 4984 99176 4984 0 _288_
rlabel metal2 99344 11256 99344 11256 0 _289_
rlabel metal2 99568 8232 99568 8232 0 _290_
rlabel metal3 60256 8008 60256 8008 0 _291_
rlabel metal2 95592 8120 95592 8120 0 _292_
rlabel metal2 62216 10192 62216 10192 0 _293_
rlabel metal3 97776 8232 97776 8232 0 _294_
rlabel metal3 100744 8120 100744 8120 0 _295_
rlabel metal2 101976 7392 101976 7392 0 _296_
rlabel metal2 97608 9408 97608 9408 0 _297_
rlabel metal2 63448 13552 63448 13552 0 _298_
rlabel metal2 95928 8512 95928 8512 0 _299_
rlabel metal2 99736 8904 99736 8904 0 _300_
rlabel metal2 102984 9464 102984 9464 0 _301_
rlabel metal2 100240 9016 100240 9016 0 _302_
rlabel metal3 44184 9016 44184 9016 0 _303_
rlabel metal2 37576 4928 37576 4928 0 _304_
rlabel metal2 63448 6160 63448 6160 0 _305_
rlabel metal2 62664 5936 62664 5936 0 _306_
rlabel metal2 23240 6384 23240 6384 0 _307_
rlabel metal2 22624 6552 22624 6552 0 _308_
rlabel metal2 12936 5040 12936 5040 0 _309_
rlabel metal2 16968 4256 16968 4256 0 _310_
rlabel metal2 19656 7504 19656 7504 0 _311_
rlabel metal2 21560 4200 21560 4200 0 _312_
rlabel metal2 27496 3472 27496 3472 0 _313_
rlabel metal2 26712 5600 26712 5600 0 _314_
rlabel metal3 38752 6104 38752 6104 0 _315_
rlabel metal2 26376 4032 26376 4032 0 _316_
rlabel metal2 27496 7504 27496 7504 0 _317_
rlabel metal3 35448 5768 35448 5768 0 _318_
rlabel metal2 30352 3752 30352 3752 0 _319_
rlabel metal2 38920 8176 38920 8176 0 _320_
rlabel metal3 32984 9016 32984 9016 0 _321_
rlabel metal3 33880 7560 33880 7560 0 _322_
rlabel metal2 45304 5824 45304 5824 0 _323_
rlabel metal2 44632 6104 44632 6104 0 _324_
rlabel metal2 47768 6608 47768 6608 0 _325_
rlabel metal3 53312 8232 53312 8232 0 _326_
rlabel metal2 37856 8344 37856 8344 0 _327_
rlabel metal2 39592 7784 39592 7784 0 _328_
rlabel metal3 49112 7336 49112 7336 0 _329_
rlabel metal2 42504 7056 42504 7056 0 _330_
rlabel metal2 44632 9464 44632 9464 0 _331_
rlabel metal2 50792 7112 50792 7112 0 _332_
rlabel metal2 47656 9240 47656 9240 0 _333_
rlabel metal2 46312 5600 46312 5600 0 _334_
rlabel metal2 51912 8316 51912 8316 0 _335_
rlabel metal2 55272 8736 55272 8736 0 _336_
rlabel metal2 54376 10640 54376 10640 0 _337_
rlabel metal2 45864 7560 45864 7560 0 _338_
rlabel metal3 57120 5992 57120 5992 0 _339_
rlabel metal2 56560 6104 56560 6104 0 _340_
rlabel metal2 57904 9240 57904 9240 0 _341_
rlabel metal2 60200 10864 60200 10864 0 _342_
rlabel metal3 60928 5992 60928 5992 0 _343_
rlabel metal3 63560 8904 63560 8904 0 _344_
rlabel metal2 63784 6608 63784 6608 0 _345_
rlabel metal2 53928 5880 53928 5880 0 clknet_0_wb_clk_i
rlabel metal2 29176 4256 29176 4256 0 clknet_3_0__leaf_wb_clk_i
rlabel metal3 22008 7336 22008 7336 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 30744 9688 30744 9688 0 clknet_3_2__leaf_wb_clk_i
rlabel metal3 51632 7896 51632 7896 0 clknet_3_3__leaf_wb_clk_i
rlabel metal2 73528 9744 73528 9744 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 73864 7616 73864 7616 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 68824 10192 68824 10192 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 73864 10192 73864 10192 0 clknet_3_7__leaf_wb_clk_i
rlabel metal3 3192 116536 3192 116536 0 io_oeb[0]
rlabel metal2 50904 116872 50904 116872 0 io_oeb[10]
rlabel metal2 54712 118146 54712 118146 0 io_oeb[11]
rlabel metal2 60312 115696 60312 115696 0 io_oeb[12]
rlabel metal2 65016 115024 65016 115024 0 io_oeb[13]
rlabel metal2 69272 117040 69272 117040 0 io_oeb[14]
rlabel metal3 73976 116536 73976 116536 0 io_oeb[15]
rlabel metal2 78232 117978 78232 117978 0 io_oeb[16]
rlabel metal2 83832 115696 83832 115696 0 io_oeb[17]
rlabel metal2 87808 115528 87808 115528 0 io_oeb[18]
rlabel metal2 93240 116592 93240 116592 0 io_oeb[19]
rlabel metal2 7672 117978 7672 117978 0 io_oeb[1]
rlabel metal3 97496 116536 97496 116536 0 io_oeb[20]
rlabel metal2 101752 117978 101752 117978 0 io_oeb[21]
rlabel metal3 107408 116536 107408 116536 0 io_oeb[22]
rlabel metal2 112280 116760 112280 116760 0 io_oeb[23]
rlabel metal2 116760 116592 116760 116592 0 io_oeb[24]
rlabel metal3 121016 116536 121016 116536 0 io_oeb[25]
rlabel metal2 125272 117978 125272 117978 0 io_oeb[26]
rlabel metal3 130928 116536 130928 116536 0 io_oeb[27]
rlabel metal2 135800 116760 135800 116760 0 io_oeb[28]
rlabel metal2 140280 116592 140280 116592 0 io_oeb[29]
rlabel metal2 13272 115696 13272 115696 0 io_oeb[2]
rlabel metal2 144984 116872 144984 116872 0 io_oeb[30]
rlabel metal2 148792 117978 148792 117978 0 io_oeb[31]
rlabel metal2 155400 116760 155400 116760 0 io_oeb[32]
rlabel metal2 159320 116816 159320 116816 0 io_oeb[33]
rlabel metal2 163800 116592 163800 116592 0 io_oeb[34]
rlabel metal2 168504 116816 168504 116816 0 io_oeb[35]
rlabel metal2 172312 117978 172312 117978 0 io_oeb[36]
rlabel metal2 18648 115808 18648 115808 0 io_oeb[3]
rlabel metal2 22232 117040 22232 117040 0 io_oeb[4]
rlabel metal2 27384 116872 27384 116872 0 io_oeb[5]
rlabel metal2 31192 117978 31192 117978 0 io_oeb[6]
rlabel metal2 36792 115696 36792 115696 0 io_oeb[7]
rlabel metal2 42280 115696 42280 115696 0 io_oeb[8]
rlabel metal2 45752 117040 45752 117040 0 io_oeb[9]
rlabel metal2 5992 116760 5992 116760 0 io_out[0]
rlabel metal3 52304 116536 52304 116536 0 io_out[10]
rlabel metal3 56728 116536 56728 116536 0 io_out[11]
rlabel metal2 61432 117208 61432 117208 0 io_out[12]
rlabel metal2 66136 116592 66136 116592 0 io_out[13]
rlabel metal2 70504 116536 70504 116536 0 io_out[14]
rlabel metal3 75824 116536 75824 116536 0 io_out[15]
rlabel metal3 80248 116536 80248 116536 0 io_out[16]
rlabel metal2 84952 117208 84952 117208 0 io_out[17]
rlabel metal2 89656 117208 89656 117208 0 io_out[18]
rlabel metal3 94192 115752 94192 115752 0 io_out[19]
rlabel metal3 9688 116536 9688 116536 0 io_out[1]
rlabel metal3 99344 116536 99344 116536 0 io_out[20]
rlabel metal3 103768 116536 103768 116536 0 io_out[21]
rlabel metal3 108304 115752 108304 115752 0 io_out[22]
rlabel metal2 113624 116760 113624 116760 0 io_out[23]
rlabel metal3 117992 115752 117992 115752 0 io_out[24]
rlabel metal3 123088 116536 123088 116536 0 io_out[25]
rlabel metal3 127400 116536 127400 116536 0 io_out[26]
rlabel metal3 132104 115752 132104 115752 0 io_out[27]
rlabel metal2 137592 116760 137592 116760 0 io_out[28]
rlabel metal3 141512 115752 141512 115752 0 io_out[29]
rlabel metal2 14392 117208 14392 117208 0 io_out[2]
rlabel metal3 146608 116536 146608 116536 0 io_out[30]
rlabel metal3 150920 116536 150920 116536 0 io_out[31]
rlabel metal2 19096 117208 19096 117208 0 io_out[3]
rlabel metal2 23464 116536 23464 116536 0 io_out[4]
rlabel metal3 28784 116536 28784 116536 0 io_out[5]
rlabel metal3 33208 116536 33208 116536 0 io_out[6]
rlabel metal2 37912 117208 37912 117208 0 io_out[7]
rlabel metal2 42616 117208 42616 117208 0 io_out[8]
rlabel metal2 46984 116536 46984 116536 0 io_out[9]
rlabel metal2 118664 5264 118664 5264 0 la_data_in[32]
rlabel metal2 120792 2198 120792 2198 0 la_data_in[33]
rlabel metal2 122360 3080 122360 3080 0 la_data_in[34]
rlabel metal2 126728 4088 126728 4088 0 la_data_in[35]
rlabel metal2 128520 3864 128520 3864 0 la_data_in[36]
rlabel metal2 131544 3584 131544 3584 0 la_data_in[37]
rlabel metal2 133392 3416 133392 3416 0 la_data_in[38]
rlabel metal2 133672 7392 133672 7392 0 la_data_in[39]
rlabel metal2 138936 4816 138936 4816 0 la_data_in[40]
rlabel metal2 138040 3640 138040 3640 0 la_data_in[41]
rlabel metal2 137368 5656 137368 5656 0 la_data_in[42]
rlabel metal2 141176 5488 141176 5488 0 la_data_in[43]
rlabel metal3 140616 3416 140616 3416 0 la_data_in[44]
rlabel metal2 142184 4816 142184 4816 0 la_data_in[45]
rlabel metal2 144984 3584 144984 3584 0 la_data_in[46]
rlabel metal2 146328 4144 146328 4144 0 la_data_in[47]
rlabel metal2 148120 3584 148120 3584 0 la_data_in[48]
rlabel metal2 149128 4816 149128 4816 0 la_data_in[49]
rlabel metal2 149352 2198 149352 2198 0 la_data_in[50]
rlabel metal3 151256 4312 151256 4312 0 la_data_in[51]
rlabel metal3 153216 3528 153216 3528 0 la_data_in[52]
rlabel metal2 155848 3584 155848 3584 0 la_data_in[53]
rlabel metal2 155960 4200 155960 4200 0 la_data_in[54]
rlabel metal3 158368 3528 158368 3528 0 la_data_in[55]
rlabel metal3 160048 3528 160048 3528 0 la_data_in[56]
rlabel metal2 161112 2534 161112 2534 0 la_data_in[57]
rlabel metal3 163240 3528 163240 3528 0 la_data_in[58]
rlabel metal3 164976 3528 164976 3528 0 la_data_in[59]
rlabel metal3 166880 3528 166880 3528 0 la_data_in[60]
rlabel metal2 169512 3584 169512 3584 0 la_data_in[61]
rlabel metal3 170184 3528 170184 3528 0 la_data_in[62]
rlabel metal3 171808 3528 171808 3528 0 la_data_in[63]
rlabel metal2 65912 2086 65912 2086 0 la_data_out[0]
rlabel metal2 82712 2058 82712 2058 0 la_data_out[10]
rlabel metal3 84784 3416 84784 3416 0 la_data_out[11]
rlabel metal2 86072 854 86072 854 0 la_data_out[12]
rlabel metal2 87752 2478 87752 2478 0 la_data_out[13]
rlabel metal3 89992 3416 89992 3416 0 la_data_out[14]
rlabel metal3 92008 3416 92008 3416 0 la_data_out[15]
rlabel metal3 93744 3528 93744 3528 0 la_data_out[16]
rlabel metal3 94920 3752 94920 3752 0 la_data_out[17]
rlabel metal3 96712 3416 96712 3416 0 la_data_out[18]
rlabel metal3 98280 4200 98280 4200 0 la_data_out[19]
rlabel metal2 67592 2086 67592 2086 0 la_data_out[1]
rlabel metal3 100128 3416 100128 3416 0 la_data_out[20]
rlabel metal3 101584 3416 101584 3416 0 la_data_out[21]
rlabel metal2 102872 2030 102872 2030 0 la_data_out[22]
rlabel metal3 105504 3416 105504 3416 0 la_data_out[23]
rlabel metal3 106680 4200 106680 4200 0 la_data_out[24]
rlabel metal3 108472 3416 108472 3416 0 la_data_out[25]
rlabel metal3 109928 4200 109928 4200 0 la_data_out[26]
rlabel metal3 111608 3416 111608 3416 0 la_data_out[27]
rlabel metal3 113512 3640 113512 3640 0 la_data_out[28]
rlabel metal3 115528 3416 115528 3416 0 la_data_out[29]
rlabel metal2 69272 2478 69272 2478 0 la_data_out[2]
rlabel metal3 117152 3640 117152 3640 0 la_data_out[30]
rlabel metal3 119168 3416 119168 3416 0 la_data_out[31]
rlabel metal2 70952 2198 70952 2198 0 la_data_out[3]
rlabel metal2 72632 2198 72632 2198 0 la_data_out[4]
rlabel metal2 74312 1246 74312 1246 0 la_data_out[5]
rlabel metal3 76440 3752 76440 3752 0 la_data_out[6]
rlabel metal3 78232 3416 78232 3416 0 la_data_out[7]
rlabel metal3 79688 3752 79688 3752 0 la_data_out[8]
rlabel metal2 81032 2198 81032 2198 0 la_data_out[9]
rlabel metal2 120232 2254 120232 2254 0 la_oenb[32]
rlabel metal2 125384 4088 125384 4088 0 la_oenb[33]
rlabel metal2 126448 3528 126448 3528 0 la_oenb[34]
rlabel metal3 127176 3528 127176 3528 0 la_oenb[35]
rlabel metal2 129024 3528 129024 3528 0 la_oenb[36]
rlabel metal2 132104 3696 132104 3696 0 la_oenb[37]
rlabel metal2 133224 7280 133224 7280 0 la_oenb[38]
rlabel metal2 135464 3584 135464 3584 0 la_oenb[39]
rlabel metal2 137144 3640 137144 3640 0 la_oenb[40]
rlabel metal2 139048 5936 139048 5936 0 la_oenb[41]
rlabel metal3 140112 3528 140112 3528 0 la_oenb[42]
rlabel metal3 139664 4312 139664 4312 0 la_oenb[43]
rlabel metal2 143304 3640 143304 3640 0 la_oenb[44]
rlabel metal3 143192 3528 143192 3528 0 la_oenb[45]
rlabel metal3 144872 3416 144872 3416 0 la_oenb[46]
rlabel metal3 146328 3528 146328 3528 0 la_oenb[47]
rlabel metal2 147112 2086 147112 2086 0 la_oenb[48]
rlabel metal2 148792 1302 148792 1302 0 la_oenb[49]
rlabel metal3 151200 3528 151200 3528 0 la_oenb[50]
rlabel metal3 152544 3416 152544 3416 0 la_oenb[51]
rlabel metal3 154504 3416 154504 3416 0 la_oenb[52]
rlabel metal3 156128 3528 156128 3528 0 la_oenb[53]
rlabel metal2 157640 3024 157640 3024 0 la_oenb[54]
rlabel metal3 159376 3416 159376 3416 0 la_oenb[55]
rlabel metal2 161672 4200 161672 4200 0 la_oenb[56]
rlabel metal3 162568 3416 162568 3416 0 la_oenb[57]
rlabel metal3 164304 3416 164304 3416 0 la_oenb[58]
rlabel metal3 166264 3416 166264 3416 0 la_oenb[59]
rlabel metal3 167944 3416 167944 3416 0 la_oenb[60]
rlabel metal2 169400 2856 169400 2856 0 la_oenb[61]
rlabel metal3 171136 3416 171136 3416 0 la_oenb[62]
rlabel metal2 172312 2086 172312 2086 0 la_oenb[63]
rlabel metal2 67648 6104 67648 6104 0 net1
rlabel metal3 88228 1064 88228 1064 0 net10
rlabel metal3 14224 5992 14224 5992 0 net100
rlabel metal2 16408 6104 16408 6104 0 net101
rlabel metal2 16072 4928 16072 4928 0 net102
rlabel metal2 8456 5600 8456 5600 0 net103
rlabel metal2 14056 5432 14056 5432 0 net104
rlabel metal2 4424 116144 4424 116144 0 net105
rlabel metal2 50008 116144 50008 116144 0 net106
rlabel metal2 54712 116144 54712 116144 0 net107
rlabel metal2 59080 115696 59080 115696 0 net108
rlabel metal2 64120 115304 64120 115304 0 net109
rlabel metal3 111328 15176 111328 15176 0 net11
rlabel metal2 68824 116144 68824 116144 0 net110
rlabel metal2 73752 116144 73752 116144 0 net111
rlabel metal2 78232 116144 78232 116144 0 net112
rlabel metal2 82600 115696 82600 115696 0 net113
rlabel metal2 87304 115192 87304 115192 0 net114
rlabel metal2 92344 116144 92344 116144 0 net115
rlabel metal2 7616 115864 7616 115864 0 net116
rlabel metal2 97272 116144 97272 116144 0 net117
rlabel metal2 101752 116144 101752 116144 0 net118
rlabel metal2 106344 116144 106344 116144 0 net119
rlabel metal2 140728 2072 140728 2072 0 net12
rlabel metal2 111160 116144 111160 116144 0 net120
rlabel metal2 115864 116144 115864 116144 0 net121
rlabel metal2 121072 115864 121072 115864 0 net122
rlabel metal2 125216 115864 125216 115864 0 net123
rlabel metal2 129864 116144 129864 116144 0 net124
rlabel metal2 134680 116144 134680 116144 0 net125
rlabel metal2 139384 116144 139384 116144 0 net126
rlabel metal2 12040 115696 12040 115696 0 net127
rlabel metal2 144088 116144 144088 116144 0 net128
rlabel metal2 148792 116144 148792 116144 0 net129
rlabel metal2 141736 3360 141736 3360 0 net13
rlabel metal2 153496 116144 153496 116144 0 net130
rlabel metal2 158200 116144 158200 116144 0 net131
rlabel metal2 162904 116144 162904 116144 0 net132
rlabel metal2 167608 116144 167608 116144 0 net133
rlabel metal2 170968 116144 170968 116144 0 net134
rlabel metal2 16968 115696 16968 115696 0 net135
rlabel metal2 21784 116144 21784 116144 0 net136
rlabel metal2 26488 116144 26488 116144 0 net137
rlabel metal2 31192 116144 31192 116144 0 net138
rlabel metal2 35560 115696 35560 115696 0 net139
rlabel metal2 141848 9408 141848 9408 0 net14
rlabel metal2 40600 115696 40600 115696 0 net140
rlabel metal2 45304 116144 45304 116144 0 net141
rlabel metal2 6776 115976 6776 115976 0 net142
rlabel metal3 53256 23576 53256 23576 0 net143
rlabel metal2 30800 3752 30800 3752 0 net144
rlabel metal2 62664 116424 62664 116424 0 net145
rlabel metal3 68768 116200 68768 116200 0 net146
rlabel metal3 69664 27384 69664 27384 0 net147
rlabel metal2 78680 116424 78680 116424 0 net148
rlabel metal3 59864 23016 59864 23016 0 net149
rlabel metal2 144592 3304 144592 3304 0 net15
rlabel metal2 90888 70840 90888 70840 0 net150
rlabel metal2 90664 116312 90664 116312 0 net151
rlabel metal3 97944 27272 97944 27272 0 net152
rlabel metal3 12040 116200 12040 116200 0 net153
rlabel metal2 50456 6944 50456 6944 0 net154
rlabel metal2 48720 10808 48720 10808 0 net155
rlabel metal2 109648 115528 109648 115528 0 net156
rlabel metal2 114408 115976 114408 115976 0 net157
rlabel metal2 117656 115584 117656 115584 0 net158
rlabel metal3 120792 116200 120792 116200 0 net159
rlabel metal2 146048 4536 146048 4536 0 net16
rlabel metal2 126952 116144 126952 116144 0 net160
rlabel metal2 131544 115528 131544 115528 0 net161
rlabel metal3 106176 1400 106176 1400 0 net162
rlabel metal2 141176 115584 141176 115584 0 net163
rlabel metal2 68152 6608 68152 6608 0 net164
rlabel metal3 146496 116424 146496 116424 0 net165
rlabel metal2 150472 116144 150472 116144 0 net166
rlabel metal2 67368 11704 67368 11704 0 net167
rlabel metal2 24808 3752 24808 3752 0 net168
rlabel metal2 24248 7224 24248 7224 0 net169
rlabel metal2 147784 2296 147784 2296 0 net17
rlabel metal2 26992 6440 26992 6440 0 net170
rlabel metal2 73080 64288 73080 64288 0 net171
rlabel metal2 27832 7896 27832 7896 0 net172
rlabel metal2 29176 6888 29176 6888 0 net173
rlabel metal2 63560 4088 63560 4088 0 net174
rlabel metal2 82152 4200 82152 4200 0 net175
rlabel metal3 83328 4424 83328 4424 0 net176
rlabel metal2 86744 3976 86744 3976 0 net177
rlabel metal2 88368 8008 88368 8008 0 net178
rlabel metal2 88144 5992 88144 5992 0 net179
rlabel metal2 148904 7000 148904 7000 0 net18
rlabel metal2 92120 3976 92120 3976 0 net180
rlabel metal2 93576 4200 93576 4200 0 net181
rlabel metal2 94472 4592 94472 4592 0 net182
rlabel metal3 95928 4872 95928 4872 0 net183
rlabel metal2 98280 5376 98280 5376 0 net184
rlabel metal2 65576 3416 65576 3416 0 net185
rlabel metal2 99904 5992 99904 5992 0 net186
rlabel metal2 102928 3528 102928 3528 0 net187
rlabel metal2 104776 3584 104776 3584 0 net188
rlabel metal2 104440 4200 104440 4200 0 net189
rlabel metal2 150808 3136 150808 3136 0 net19
rlabel metal2 104440 5488 104440 5488 0 net190
rlabel metal2 108248 4760 108248 4760 0 net191
rlabel metal2 110656 6440 110656 6440 0 net192
rlabel metal2 112840 4032 112840 4032 0 net193
rlabel metal2 112392 3976 112392 3976 0 net194
rlabel metal2 115192 7616 115192 7616 0 net195
rlabel metal3 64680 4368 64680 4368 0 net196
rlabel metal2 115752 8736 115752 8736 0 net197
rlabel metal3 118440 9128 118440 9128 0 net198
rlabel metal2 67760 8008 67760 8008 0 net199
rlabel metal3 68768 13608 68768 13608 0 net2
rlabel metal2 151312 4536 151312 4536 0 net20
rlabel metal2 73808 3528 73808 3528 0 net200
rlabel metal2 74312 5544 74312 5544 0 net201
rlabel metal2 75656 4368 75656 4368 0 net202
rlabel metal2 77784 8008 77784 8008 0 net203
rlabel metal2 79184 5992 79184 5992 0 net204
rlabel metal2 80248 6832 80248 6832 0 net205
rlabel metal2 6888 4144 6888 4144 0 net206
rlabel metal2 11256 5656 11256 5656 0 net207
rlabel metal2 30968 6160 30968 6160 0 net208
rlabel metal2 32088 3808 32088 3808 0 net209
rlabel metal2 153496 2240 153496 2240 0 net21
rlabel metal2 34440 5544 34440 5544 0 net210
rlabel metal2 34328 6216 34328 6216 0 net211
rlabel metal2 43736 7896 43736 7896 0 net212
rlabel metal2 49112 4536 49112 4536 0 net213
rlabel metal2 40264 5964 40264 5964 0 net214
rlabel metal2 40824 7224 40824 7224 0 net215
rlabel metal3 45304 6552 45304 6552 0 net216
rlabel metal2 44968 5320 44968 5320 0 net217
rlabel metal2 11704 3080 11704 3080 0 net218
rlabel metal2 49672 6496 49672 6496 0 net219
rlabel metal2 155624 2408 155624 2408 0 net22
rlabel metal2 48104 5264 48104 5264 0 net220
rlabel metal2 45528 3864 45528 3864 0 net221
rlabel metal2 51464 5936 51464 5936 0 net222
rlabel metal2 54152 4760 54152 4760 0 net223
rlabel metal2 56784 5208 56784 5208 0 net224
rlabel metal2 55720 4760 55720 4760 0 net225
rlabel metal2 57960 3976 57960 3976 0 net226
rlabel metal2 59864 5964 59864 5964 0 net227
rlabel metal3 60648 6440 60648 6440 0 net228
rlabel metal2 14952 4592 14952 4592 0 net229
rlabel metal2 156296 7504 156296 7504 0 net23
rlabel metal2 63448 3528 63448 3528 0 net230
rlabel metal2 65128 6104 65128 6104 0 net231
rlabel metal2 18984 4368 18984 4368 0 net232
rlabel metal2 20776 5824 20776 5824 0 net233
rlabel metal2 22456 3472 22456 3472 0 net234
rlabel metal3 25536 4424 25536 4424 0 net235
rlabel metal2 23800 4760 23800 4760 0 net236
rlabel metal3 25928 3528 25928 3528 0 net237
rlabel metal2 28672 6552 28672 6552 0 net238
rlabel metal2 177128 116312 177128 116312 0 net239
rlabel metal2 158648 2352 158648 2352 0 net24
rlabel metal2 155176 115864 155176 115864 0 net240
rlabel metal2 160440 116648 160440 116648 0 net241
rlabel metal3 164696 116312 164696 116312 0 net242
rlabel metal3 169792 116312 169792 116312 0 net243
rlabel metal2 174328 117096 174328 117096 0 net244
rlabel metal3 178360 115864 178360 115864 0 net245
rlabel metal2 172872 2590 172872 2590 0 net246
rlabel metal2 173432 1246 173432 1246 0 net247
rlabel metal2 173992 2030 173992 2030 0 net248
rlabel metal2 119672 2030 119672 2030 0 net249
rlabel metal2 160440 7056 160440 7056 0 net25
rlabel metal2 121352 1582 121352 1582 0 net250
rlabel metal2 123032 1134 123032 1134 0 net251
rlabel metal2 124824 5992 124824 5992 0 net252
rlabel metal2 126392 1582 126392 1582 0 net253
rlabel metal3 128968 3864 128968 3864 0 net254
rlabel metal2 129752 2058 129752 2058 0 net255
rlabel metal2 131544 5208 131544 5208 0 net256
rlabel metal2 133112 2198 133112 2198 0 net257
rlabel metal2 134792 2030 134792 2030 0 net258
rlabel metal2 136472 3598 136472 3598 0 net259
rlabel metal2 161336 9072 161336 9072 0 net26
rlabel metal2 138152 854 138152 854 0 net260
rlabel metal2 139832 1582 139832 1582 0 net261
rlabel metal2 141512 1862 141512 1862 0 net262
rlabel metal2 143192 3374 143192 3374 0 net263
rlabel metal2 144872 3598 144872 3598 0 net264
rlabel metal2 146552 3374 146552 3374 0 net265
rlabel metal2 148232 2310 148232 2310 0 net266
rlabel metal2 149912 1582 149912 1582 0 net267
rlabel metal2 151592 1582 151592 1582 0 net268
rlabel metal2 153272 2590 153272 2590 0 net269
rlabel metal2 163464 10920 163464 10920 0 net27
rlabel metal2 154952 2590 154952 2590 0 net270
rlabel metal2 156632 2086 156632 2086 0 net271
rlabel metal2 158312 1414 158312 1414 0 net272
rlabel metal2 159992 2590 159992 2590 0 net273
rlabel metal2 161672 1470 161672 1470 0 net274
rlabel metal2 163352 1078 163352 1078 0 net275
rlabel metal2 165032 2590 165032 2590 0 net276
rlabel metal2 166712 2590 166712 2590 0 net277
rlabel metal2 168392 1526 168392 1526 0 net278
rlabel metal2 170072 2590 170072 2590 0 net279
rlabel metal2 159208 3752 159208 3752 0 net28
rlabel metal2 171752 2590 171752 2590 0 net280
rlabel metal2 167384 12096 167384 12096 0 net29
rlabel metal4 70280 8736 70280 8736 0 net3
rlabel metal2 169232 3304 169232 3304 0 net30
rlabel metal2 170408 7616 170408 7616 0 net31
rlabel metal2 172200 6832 172200 6832 0 net32
rlabel metal3 122248 4872 122248 4872 0 net33
rlabel metal2 125160 3248 125160 3248 0 net34
rlabel metal3 125832 3304 125832 3304 0 net35
rlabel metal3 128856 3752 128856 3752 0 net36
rlabel metal2 143360 4312 143360 4312 0 net37
rlabel metal2 132440 3808 132440 3808 0 net38
rlabel metal2 133560 4368 133560 4368 0 net39
rlabel metal3 69776 13048 69776 13048 0 net4
rlabel metal3 134792 4984 134792 4984 0 net40
rlabel metal3 134400 3304 134400 3304 0 net41
rlabel metal2 139496 3304 139496 3304 0 net42
rlabel metal2 139944 3192 139944 3192 0 net43
rlabel metal2 140392 3864 140392 3864 0 net44
rlabel metal3 142240 3304 142240 3304 0 net45
rlabel metal2 143864 3080 143864 3080 0 net46
rlabel metal2 145208 4480 145208 4480 0 net47
rlabel metal3 145432 3304 145432 3304 0 net48
rlabel metal2 138152 6160 138152 6160 0 net49
rlabel metal3 71568 4312 71568 4312 0 net5
rlabel metal3 148904 4424 148904 4424 0 net50
rlabel metal3 147336 4256 147336 4256 0 net51
rlabel metal2 140112 7336 140112 7336 0 net52
rlabel metal2 148008 4088 148008 4088 0 net53
rlabel metal2 156520 3584 156520 3584 0 net54
rlabel metal3 150808 4368 150808 4368 0 net55
rlabel metal2 146104 5712 146104 5712 0 net56
rlabel metal2 161392 3304 161392 3304 0 net57
rlabel metal2 162568 2800 162568 2800 0 net58
rlabel metal2 164360 5432 164360 5432 0 net59
rlabel metal2 131208 2912 131208 2912 0 net6
rlabel metal2 139720 3304 139720 3304 0 net60
rlabel metal2 168280 3024 168280 3024 0 net61
rlabel metal2 169064 3024 169064 3024 0 net62
rlabel metal2 171304 5656 171304 5656 0 net63
rlabel metal2 144984 4592 144984 4592 0 net64
rlabel metal2 8344 2296 8344 2296 0 net65
rlabel metal2 7896 5040 7896 5040 0 net66
rlabel metal3 21196 4536 21196 4536 0 net67
rlabel metal2 29960 9352 29960 9352 0 net68
rlabel metal2 28504 8512 28504 8512 0 net69
rlabel metal2 63672 4480 63672 4480 0 net7
rlabel metal2 29736 9688 29736 9688 0 net70
rlabel metal2 32928 6104 32928 6104 0 net71
rlabel metal2 36792 4200 36792 4200 0 net72
rlabel metal2 37968 7672 37968 7672 0 net73
rlabel metal2 39144 4704 39144 4704 0 net74
rlabel metal2 120792 23548 120792 23548 0 net75
rlabel metal2 40992 6552 40992 6552 0 net76
rlabel metal2 52136 4816 52136 4816 0 net77
rlabel metal3 20160 3696 20160 3696 0 net78
rlabel metal2 46816 9576 46816 9576 0 net79
rlabel metal2 133896 3752 133896 3752 0 net8
rlabel metal3 47936 9240 47936 9240 0 net80
rlabel metal2 47376 7672 47376 7672 0 net81
rlabel metal2 44744 13944 44744 13944 0 net82
rlabel metal2 46760 6104 46760 6104 0 net83
rlabel metal2 49280 4984 49280 4984 0 net84
rlabel metal2 55776 7672 55776 7672 0 net85
rlabel metal3 57344 6552 57344 6552 0 net86
rlabel metal2 57792 8120 57792 8120 0 net87
rlabel metal2 60760 3752 60760 3752 0 net88
rlabel metal3 26040 6384 26040 6384 0 net89
rlabel metal2 136024 2856 136024 2856 0 net9
rlabel metal2 58016 4536 58016 4536 0 net90
rlabel metal2 65352 7056 65352 7056 0 net91
rlabel metal2 40488 6776 40488 6776 0 net92
rlabel metal3 71176 10584 71176 10584 0 net93
rlabel metal2 21784 3584 21784 3584 0 net94
rlabel metal2 73360 4312 73360 4312 0 net95
rlabel metal2 24472 9464 24472 9464 0 net96
rlabel metal2 23128 11592 23128 11592 0 net97
rlabel metal2 25648 3304 25648 3304 0 net98
rlabel metal3 24696 6048 24696 6048 0 net99
rlabel metal2 5992 4606 5992 4606 0 wb_clk_i
rlabel metal2 6552 2142 6552 2142 0 wb_rst_i
rlabel metal2 7112 2478 7112 2478 0 wbs_ack_o
rlabel metal2 7672 2926 7672 2926 0 wbs_cyc_i
rlabel metal2 10024 4312 10024 4312 0 wbs_dat_i[0]
rlabel metal2 29568 6552 29568 6552 0 wbs_dat_i[10]
rlabel metal3 29456 3528 29456 3528 0 wbs_dat_i[11]
rlabel metal2 29512 3640 29512 3640 0 wbs_dat_i[12]
rlabel metal2 31528 6608 31528 6608 0 wbs_dat_i[13]
rlabel metal2 31752 5712 31752 5712 0 wbs_dat_i[14]
rlabel metal2 37464 7448 37464 7448 0 wbs_dat_i[15]
rlabel metal2 38920 5656 38920 5656 0 wbs_dat_i[16]
rlabel metal3 40040 6552 40040 6552 0 wbs_dat_i[17]
rlabel metal3 41384 6552 41384 6552 0 wbs_dat_i[18]
rlabel metal2 44856 7896 44856 7896 0 wbs_dat_i[19]
rlabel metal2 11256 3864 11256 3864 0 wbs_dat_i[1]
rlabel metal2 46424 8064 46424 8064 0 wbs_dat_i[20]
rlabel metal2 47432 2478 47432 2478 0 wbs_dat_i[21]
rlabel metal3 47880 7448 47880 7448 0 wbs_dat_i[22]
rlabel metal2 44408 4592 44408 4592 0 wbs_dat_i[23]
rlabel metal2 46648 5768 46648 5768 0 wbs_dat_i[24]
rlabel metal3 51464 4984 51464 4984 0 wbs_dat_i[25]
rlabel metal2 55832 4102 55832 4102 0 wbs_dat_i[26]
rlabel metal2 57680 6552 57680 6552 0 wbs_dat_i[27]
rlabel metal2 57512 7896 57512 7896 0 wbs_dat_i[28]
rlabel metal2 60424 5488 60424 5488 0 wbs_dat_i[29]
rlabel metal2 14168 5376 14168 5376 0 wbs_dat_i[2]
rlabel metal3 60032 4312 60032 4312 0 wbs_dat_i[30]
rlabel metal2 65016 4368 65016 4368 0 wbs_dat_i[31]
rlabel metal3 15456 3528 15456 3528 0 wbs_dat_i[3]
rlabel metal2 18480 4312 18480 4312 0 wbs_dat_i[4]
rlabel metal2 20552 3262 20552 3262 0 wbs_dat_i[5]
rlabel metal2 22456 4928 22456 4928 0 wbs_dat_i[6]
rlabel metal2 24080 5880 24080 5880 0 wbs_dat_i[7]
rlabel metal3 24136 4312 24136 4312 0 wbs_dat_i[8]
rlabel metal2 25480 3640 25480 3640 0 wbs_dat_i[9]
rlabel metal2 10472 2198 10472 2198 0 wbs_dat_o[0]
rlabel metal2 29512 854 29512 854 0 wbs_dat_o[10]
rlabel metal2 31192 2982 31192 2982 0 wbs_dat_o[11]
rlabel metal2 32872 2086 32872 2086 0 wbs_dat_o[12]
rlabel metal2 34552 2478 34552 2478 0 wbs_dat_o[13]
rlabel metal2 36232 2086 36232 2086 0 wbs_dat_o[14]
rlabel metal2 37912 2198 37912 2198 0 wbs_dat_o[15]
rlabel metal2 39592 2198 39592 2198 0 wbs_dat_o[16]
rlabel metal2 41272 2198 41272 2198 0 wbs_dat_o[17]
rlabel metal2 42952 854 42952 854 0 wbs_dat_o[18]
rlabel metal2 44632 1470 44632 1470 0 wbs_dat_o[19]
rlabel metal2 12712 2198 12712 2198 0 wbs_dat_o[1]
rlabel metal2 46312 2030 46312 2030 0 wbs_dat_o[20]
rlabel metal2 47992 1246 47992 1246 0 wbs_dat_o[21]
rlabel metal2 49672 2086 49672 2086 0 wbs_dat_o[22]
rlabel metal2 51352 3654 51352 3654 0 wbs_dat_o[23]
rlabel metal2 53032 2198 53032 2198 0 wbs_dat_o[24]
rlabel metal2 54712 2478 54712 2478 0 wbs_dat_o[25]
rlabel metal2 56392 2086 56392 2086 0 wbs_dat_o[26]
rlabel metal2 58072 2086 58072 2086 0 wbs_dat_o[27]
rlabel metal2 59752 2086 59752 2086 0 wbs_dat_o[28]
rlabel metal2 61432 2198 61432 2198 0 wbs_dat_o[29]
rlabel metal2 14952 2086 14952 2086 0 wbs_dat_o[2]
rlabel metal2 63112 2198 63112 2198 0 wbs_dat_o[30]
rlabel metal2 64792 1414 64792 1414 0 wbs_dat_o[31]
rlabel metal2 17192 2086 17192 2086 0 wbs_dat_o[3]
rlabel metal2 19432 2982 19432 2982 0 wbs_dat_o[4]
rlabel metal2 21112 2086 21112 2086 0 wbs_dat_o[5]
rlabel metal2 22792 1638 22792 1638 0 wbs_dat_o[6]
rlabel metal2 24472 2478 24472 2478 0 wbs_dat_o[7]
rlabel metal2 26152 2086 26152 2086 0 wbs_dat_o[8]
rlabel metal2 27832 2982 27832 2982 0 wbs_dat_o[9]
rlabel metal2 10808 4704 10808 4704 0 wbs_sel_i[0]
rlabel metal2 13272 3318 13272 3318 0 wbs_sel_i[1]
rlabel metal2 15624 5880 15624 5880 0 wbs_sel_i[2]
rlabel metal2 15848 4144 15848 4144 0 wbs_sel_i[3]
rlabel metal2 8120 5768 8120 5768 0 wbs_stb_i
rlabel metal2 9576 4256 9576 4256 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 180000 120000
<< end >>
