magic
tech gf180mcuC
magscale 1 5
timestamp 1670117523
<< obsm1 >>
rect 672 1538 89320 58505
<< metal2 >>
rect 1568 59600 1624 60000
rect 4368 59600 4424 60000
rect 7168 59600 7224 60000
rect 9968 59600 10024 60000
rect 12768 59600 12824 60000
rect 15568 59600 15624 60000
rect 18368 59600 18424 60000
rect 21168 59600 21224 60000
rect 23968 59600 24024 60000
rect 26768 59600 26824 60000
rect 29568 59600 29624 60000
rect 32368 59600 32424 60000
rect 35168 59600 35224 60000
rect 37968 59600 38024 60000
rect 40768 59600 40824 60000
rect 43568 59600 43624 60000
rect 46368 59600 46424 60000
rect 49168 59600 49224 60000
rect 51968 59600 52024 60000
rect 54768 59600 54824 60000
rect 57568 59600 57624 60000
rect 60368 59600 60424 60000
rect 63168 59600 63224 60000
rect 65968 59600 66024 60000
rect 68768 59600 68824 60000
rect 71568 59600 71624 60000
rect 74368 59600 74424 60000
rect 77168 59600 77224 60000
rect 79968 59600 80024 60000
rect 82768 59600 82824 60000
rect 85568 59600 85624 60000
rect 88368 59600 88424 60000
rect 4648 0 4704 400
rect 13608 0 13664 400
rect 22568 0 22624 400
rect 31528 0 31584 400
rect 40488 0 40544 400
rect 49448 0 49504 400
rect 58408 0 58464 400
rect 67368 0 67424 400
rect 76328 0 76384 400
rect 85288 0 85344 400
<< obsm2 >>
rect 1654 59570 4338 59600
rect 4454 59570 7138 59600
rect 7254 59570 9938 59600
rect 10054 59570 12738 59600
rect 12854 59570 15538 59600
rect 15654 59570 18338 59600
rect 18454 59570 21138 59600
rect 21254 59570 23938 59600
rect 24054 59570 26738 59600
rect 26854 59570 29538 59600
rect 29654 59570 32338 59600
rect 32454 59570 35138 59600
rect 35254 59570 37938 59600
rect 38054 59570 40738 59600
rect 40854 59570 43538 59600
rect 43654 59570 46338 59600
rect 46454 59570 49138 59600
rect 49254 59570 51938 59600
rect 52054 59570 54738 59600
rect 54854 59570 57538 59600
rect 57654 59570 60338 59600
rect 60454 59570 63138 59600
rect 63254 59570 65938 59600
rect 66054 59570 68738 59600
rect 68854 59570 71538 59600
rect 71654 59570 74338 59600
rect 74454 59570 77138 59600
rect 77254 59570 79938 59600
rect 80054 59570 82738 59600
rect 82854 59570 85538 59600
rect 85654 59570 88338 59600
rect 88454 59570 88466 59600
rect 1582 430 88466 59570
rect 1582 400 4618 430
rect 4734 400 13578 430
rect 13694 400 22538 430
rect 22654 400 31498 430
rect 31614 400 40458 430
rect 40574 400 49418 430
rect 49534 400 58378 430
rect 58494 400 67338 430
rect 67454 400 76298 430
rect 76414 400 85258 430
rect 85374 400 88466 430
<< obsm3 >>
rect 2233 1414 88135 58506
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
rect 86704 1538 86864 58438
<< obsm4 >>
rect 36974 4153 40594 56327
rect 40814 4153 40866 56327
<< labels >>
rlabel metal2 s 76328 0 76384 400 6 clk
port 1 nsew signal input
rlabel metal2 s 1568 59600 1624 60000 6 fn[0]
port 2 nsew signal output
rlabel metal2 s 29568 59600 29624 60000 6 fn[10]
port 3 nsew signal output
rlabel metal2 s 32368 59600 32424 60000 6 fn[11]
port 4 nsew signal output
rlabel metal2 s 35168 59600 35224 60000 6 fn[12]
port 5 nsew signal output
rlabel metal2 s 37968 59600 38024 60000 6 fn[13]
port 6 nsew signal output
rlabel metal2 s 40768 59600 40824 60000 6 fn[14]
port 7 nsew signal output
rlabel metal2 s 43568 59600 43624 60000 6 fn[15]
port 8 nsew signal output
rlabel metal2 s 46368 59600 46424 60000 6 fn[16]
port 9 nsew signal output
rlabel metal2 s 49168 59600 49224 60000 6 fn[17]
port 10 nsew signal output
rlabel metal2 s 51968 59600 52024 60000 6 fn[18]
port 11 nsew signal output
rlabel metal2 s 54768 59600 54824 60000 6 fn[19]
port 12 nsew signal output
rlabel metal2 s 4368 59600 4424 60000 6 fn[1]
port 13 nsew signal output
rlabel metal2 s 57568 59600 57624 60000 6 fn[20]
port 14 nsew signal output
rlabel metal2 s 60368 59600 60424 60000 6 fn[21]
port 15 nsew signal output
rlabel metal2 s 63168 59600 63224 60000 6 fn[22]
port 16 nsew signal output
rlabel metal2 s 65968 59600 66024 60000 6 fn[23]
port 17 nsew signal output
rlabel metal2 s 68768 59600 68824 60000 6 fn[24]
port 18 nsew signal output
rlabel metal2 s 71568 59600 71624 60000 6 fn[25]
port 19 nsew signal output
rlabel metal2 s 74368 59600 74424 60000 6 fn[26]
port 20 nsew signal output
rlabel metal2 s 77168 59600 77224 60000 6 fn[27]
port 21 nsew signal output
rlabel metal2 s 79968 59600 80024 60000 6 fn[28]
port 22 nsew signal output
rlabel metal2 s 82768 59600 82824 60000 6 fn[29]
port 23 nsew signal output
rlabel metal2 s 7168 59600 7224 60000 6 fn[2]
port 24 nsew signal output
rlabel metal2 s 85568 59600 85624 60000 6 fn[30]
port 25 nsew signal output
rlabel metal2 s 88368 59600 88424 60000 6 fn[31]
port 26 nsew signal output
rlabel metal2 s 9968 59600 10024 60000 6 fn[3]
port 27 nsew signal output
rlabel metal2 s 12768 59600 12824 60000 6 fn[4]
port 28 nsew signal output
rlabel metal2 s 15568 59600 15624 60000 6 fn[5]
port 29 nsew signal output
rlabel metal2 s 18368 59600 18424 60000 6 fn[6]
port 30 nsew signal output
rlabel metal2 s 21168 59600 21224 60000 6 fn[7]
port 31 nsew signal output
rlabel metal2 s 23968 59600 24024 60000 6 fn[8]
port 32 nsew signal output
rlabel metal2 s 26768 59600 26824 60000 6 fn[9]
port 33 nsew signal output
rlabel metal2 s 4648 0 4704 400 6 n[0]
port 34 nsew signal input
rlabel metal2 s 13608 0 13664 400 6 n[1]
port 35 nsew signal input
rlabel metal2 s 22568 0 22624 400 6 n[2]
port 36 nsew signal input
rlabel metal2 s 31528 0 31584 400 6 n[3]
port 37 nsew signal input
rlabel metal2 s 40488 0 40544 400 6 n[4]
port 38 nsew signal input
rlabel metal2 s 49448 0 49504 400 6 n[5]
port 39 nsew signal input
rlabel metal2 s 58408 0 58464 400 6 n[6]
port 40 nsew signal input
rlabel metal2 s 67368 0 67424 400 6 n[7]
port 41 nsew signal input
rlabel metal2 s 85288 0 85344 400 6 st
port 42 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 44 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 44 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 44 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 44 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vss
port 44 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 58438 6 vss
port 44 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2916130
string GDS_FILE /home/ivan/Documentos/global_foundries/gf180-demo/caravel_user_project/openlane/user_proj_example/runs/22_12_03_20_30/results/signoff/fibonacci.magic.gds
string GDS_START 253956
<< end >>

